/*TOPOLOGY*/
`define MESH_TOPOLOGY_X              5//`DSU_MAX_X_NUM
`define MESH_TOPOLOGY_Y              2//`DSU_MAX_Y_NUM

`define NOC_ROUTECOMPX_W             $clog2(`MESH_TOPOLOGY_X)
`define NOC_ROUTECOMPY_W             $clog2(`MESH_TOPOLOGY_Y)

/*DIRECTION PORTS*/
`define DIRECTION_E                  0
`define DIRECTION_W                  1
`define DIRECTION_N                  2
`define DIRECTION_S                  3
`define DEVICE_P0                    4
`define DEVICE_P1                    5
`define DEVICE_P2                    6
`define DEVICE_P3                    7

`define DEVICE_PORT_NUM              4
`define TOTAL_PORT_NUM               8
`define CROSSBAR_MUX_NUM             8

`define DLB_PORT_NUM                 8
`define DLB_CROSSBAR_MUX_NUM         8

/*CHANNEL TYPE*/
`define CHANNEL_REQ                  0
`define CHANNEL_RSP                  1
`define CHANNEL_SNP                  2
`define CHANNEL_DAT                  3
`define CHANNEL_DLB                  4

/*CRD WIDTH*/
`define ROUTER_CRD_WIDTH             4
`define DEVICE_CRD_WIDTH             15

`define MESH_REQ_FLIT_WIDTH          `DSU_CHI_REQ_FLIT_WIDTH
`define MESH_RSP_FLIT_WIDTH          `DSU_CHI_RSP_FLIT_WIDTH
`define MESH_SNP_FLIT_WIDTH          `DSU_CHI_SNP_FLIT_WIDTH
`define MESH_DAT_FLIT_WIDTH          `DSU_CHI_DAT_FLIT_WIDTH
`define MESH_DLB_FLIT_WIDTH          `DSU_DLB_FLIT_WIDTH
`define DSU_CHI_DLB_FLIT_WIDTH       `DSU_DLB_FLIT_WIDTH

`define RNFBESAM_REQ_FLIT_WIDTH      `DSU_CHI_RNFBESAM_REQ_FLIT_WIDTH
`define RNFBESAM_RSP_FLIT_WIDTH      `DSU_CHI_RNFBESAM_RSP_FLIT_WIDTH
`define RNFBESAM_SNP_FLIT_WIDTH      `DSU_CHI_RNFBESAM_SNP_FLIT_WIDTH
`define RNFBESAM_DAT_FLIT_WIDTH      `DSU_CHI_RNFBESAM_DAT_FLIT_WIDTH
`define HNDBESAM_DLB_FLIT_WIDTH      `DSU_DLB_FLIT_WIDTH

/*TGTID MACRO*/
`define NOC_ROUTE_WIDTH              `DSU_NODEID_WIDTH
`define NOC_ROUTE_DEVICEID_WIDTH     `DSU_MXP_DEVICEID_WIDTH_PARAM
`define NOC_ROUTE_PORTID_WIDTH       `DSU_MXP_PORTID_WIDTH_PARAM
`define NOC_ROUTE_YID_WIDTH          `DSU_MXP_YID_WIDTH_PARAM
`define NOC_ROUTE_XID_WIDTH          `DSU_MXP_XID_WIDTH_PARAM

`define NOC_ROUTE_DEVICEID_RIGHT     0
`define NOC_ROUTE_DEVICEID_LEFT      (`NOC_ROUTE_DEVICEID_RIGHT + `NOC_ROUTE_DEVICEID_WIDTH -1)
`define NOC_ROUTE_PORTID_RIGHT       (`NOC_ROUTE_DEVICEID_LEFT  + 1)
`define NOC_ROUTE_PORTID_LEFT        (`NOC_ROUTE_PORTID_RIGHT   + `NOC_ROUTE_PORTID_WIDTH   -1)
`define NOC_ROUTE_YID_RIGHT          (`NOC_ROUTE_PORTID_LEFT    + 1)
`define NOC_ROUTE_YID_LEFT           (`NOC_ROUTE_YID_RIGHT      + `NOC_ROUTE_YID_WIDTH      -1)
`define NOC_ROUTE_XID_RIGHT          (`NOC_ROUTE_YID_LEFT       + 1)
`define NOC_ROUTE_XID_LEFT           (`NOC_ROUTE_XID_RIGHT      + `NOC_ROUTE_XID_WIDTH      -1)

`define NOC_ROUTE_PORTID_RANGE       `NOC_ROUTE_PORTID_LEFT    : `NOC_ROUTE_PORTID_RIGHT     
`define NOC_ROUTE_YID_RANGE          `NOC_ROUTE_YID_LEFT       : `NOC_ROUTE_YID_RIGHT        
`define NOC_ROUTE_XID_RANGE          `NOC_ROUTE_XID_LEFT       : `NOC_ROUTE_XID_RIGHT        
`define NOC_ROUTE_NID_RANGE          `NOC_ROUTE_XID_LEFT       : 0

`define DLB_ROUTE_WIDTH              `DSU_DLB_MESH_TGTID_WIDTH
`define DLB_ROUTE_DEVICEID_WIDTH     `DSU_DLB_MESH_DEVICEID_WIDTH
`define DLB_ROUTE_PORTID_WIDTH       `DSU_DLB_MESH_PORTID_WIDTH
`define DLB_ROUTE_TODEV_WIDTH        `DSU_DLB_MESH_TODEV_WIDTH
`define DLB_ROUTE_YID_WIDTH          `DSU_DLB_MESH_YID_WIDTH
`define DLB_ROUTE_XID_WIDTH          `DSU_DLB_MESH_XID_WIDTH

`define DLB_ROUTE_DEVICEID_RIGHT     0
`define DLB_ROUTE_DEVICEID_LEFT      (`DLB_ROUTE_DEVICEID_RIGHT + `DLB_ROUTE_DEVICEID_WIDTH -1)
`define DLB_ROUTE_PORTID_RIGHT       (`DLB_ROUTE_DEVICEID_LEFT+1)
`define DLB_ROUTE_PORTID_LEFT        (`DLB_ROUTE_PORTID_RIGHT+`DSU_DLB_MESH_PORTID_WIDTH-1)
`define DLB_ROUTE_TODEV_RIGHT        (`DLB_ROUTE_PORTID_LEFT+1)
`define DLB_ROUTE_TODEV_LEFT         (`DLB_ROUTE_TODEV_RIGHT+`DSU_DLB_MESH_TODEV_WIDTH-1)
`define DLB_ROUTE_YID_RIGHT          (`DLB_ROUTE_TODEV_LEFT+ 1)
`define DLB_ROUTE_YID_LEFT           (`DLB_ROUTE_YID_RIGHT + `DLB_ROUTE_YID_WIDTH -1)
`define DLB_ROUTE_XID_RIGHT          (`DLB_ROUTE_YID_LEFT + 1)
`define DLB_ROUTE_XID_LEFT           (`DLB_ROUTE_XID_RIGHT + `DLB_ROUTE_XID_WIDTH -1)

`define DLB_ROUTE_DEVICEID_RANGE     `DLB_ROUTE_DEVICEID_LEFT:`DLB_ROUTE_DEVICEID_RIGHT 
`define DLB_ROUTE_PORTID_RANGE       `DLB_ROUTE_PORTID_LEFT:`DLB_ROUTE_PORTID_RIGHT
`define DLB_ROUTE_TODEV_RANGE         `DLB_ROUTE_TODEV_LEFT:`DLB_ROUTE_TODEV_RIGHT
`define DLB_ROUTE_YID_RANGE          `DLB_ROUTE_YID_LEFT:`DLB_ROUTE_YID_RIGHT    
`define DLB_ROUTE_XID_RANGE          `DLB_ROUTE_XID_LEFT:`DLB_ROUTE_XID_RIGHT     

/*REQ FLIT*/
`define CHI_REQ_PCRDRETURN_OPCODE   `DSU_CHI_REQ_OP_PCRDRETURN
// CHI B
// `define REQ_FLIT_QOS_RANGE           `DSU_CHI_REQ_FLIT_QOS_RANGE
// `define REQ_FLIT_TGTID_RANGE         `DSU_CHI_REQ_FLIT_TGTID_RANGE
// `define REQ_FLIT_SRCID_RANGE         `DSU_CHI_REQ_FLIT_SRCID_RANGE
// `define REQ_FLIT_TXNID_RANGE         `DSU_CHI_REQ_FLIT_TXNID_RANGE
// `define REQ_FLIT_RNID_RANGE          `DSU_CHI_REQ_FLIT_RNID_RANGE
// `define REQ_FLIT_STASHNIDV_RANGE     `DSU_CHI_REQ_FLIT_STASHNIDV_RANGE
// `define REQ_FLIT_RETURNTXNID_RANGE   `DSU_CHI_REQ_FLIT_RETURNTXNID_RANGE
// `define REQ_FLIT_OPCODE_RANGE        `DSU_CHI_REQ_FLIT_OPCODE_RANGE
// `define REQ_FLIT_SIZE_RANGE          `DSU_CHI_REQ_FLIT_SIZE_RANGE
// `define REQ_FLIT_ADDR_RANGE          `DSU_CHI_REQ_FLIT_ADDR_RANGE
// `define REQ_FLIT_NS_RANGE            `DSU_CHI_REQ_FLIT_NS_RANGE
// `define REQ_FLIT_LS_RANGE            `DSU_CHI_REQ_FLIT_LS_RANGE
// `define REQ_FLIT_ALLOWRETRY_RANGE    `DSU_CHI_REQ_FLIT_ALLOWRETRY_RANGE
// `define REQ_FLIT_ORDER_RANGE         `DSU_CHI_REQ_FLIT_ORDER_RANGE
// `define REQ_FLIT_PCRDTYPE_RANGE      `DSU_CHI_REQ_FLIT_PCRDTYPE_RANGE
// `define REQ_FLIT_MEMATTR_RANGE       `DSU_CHI_REQ_FLIT_MEMATTR_RANGE
// `define REQ_FLIT_SNPATTR_RANGE       `DSU_CHI_REQ_FLIT_SNPATTR_RANGE
// `define REQ_FLIT_LPID_RANGE          `DSU_CHI_REQ_FLIT_LPID_RANGE
// `define REQ_FLIT_EXCL_RANGE          `DSU_CHI_REQ_FLIT_EXCL_RANGE
// `define REQ_FLIT_EXPCOMPACK_RANGE    `DSU_CHI_REQ_FLIT_EXPCOMPACK_RANGE
// `define REQ_FLIT_TRACETAG_RANGE      `DSU_CHI_REQ_FLIT_TRACETAG_RANGE
// `define REQ_FLIT_RSVD_RANGE          `DSU_CHI_REQ_FLIT_RSVD_RANGE
// `define REQ_FLIT_SRCTYPE_RANGE       `DSU_CHI_REQ_FLIT_SRCTYPE_RANGE
// `define REQ_FLIT_LDID_RANGE          `DSU_CHI_REQ_FLIT_LDID_RANGE

//CHI E
`define REQ_FLIT_QOS_RANGE              `DSU_CHI_REQ_FLIT_QOS_RANGE    
`define REQ_FLIT_DEVICEID_RANGE         `DSU_CHI_REQ_FLIT_DEVICEID_RANGE         
`define REQ_FLIT_PORTID_RANGE           `DSU_CHI_REQ_FLIT_PORTID_RANGE       
`define REQ_FLIT_YID_RANGE              `DSU_CHI_REQ_FLIT_YID_RANGE    
`define REQ_FLIT_XID_RANGE              `DSU_CHI_REQ_FLIT_XID_RANGE    
`define REQ_FLIT_MESHID_RANGE           `DSU_CHI_REQ_FLIT_MESHID_RANGE       
`define REQ_FLIT_TGTID_RANGE            `DSU_CHI_REQ_FLIT_TGTID_RANGE      
`define REQ_FLIT_SRCID_RANGE            `DSU_CHI_REQ_FLIT_SRCID_RANGE      
`define REQ_FLIT_TXNID_RANGE            `DSU_CHI_REQ_FLIT_TXNID_RANGE      
`define REQ_FLIT_RNID_RANGE             `DSU_CHI_REQ_FLIT_RNID_RANGE     
`define REQ_FLIT_STASHNIDV_RANGE        `DSU_CHI_REQ_FLIT_STASHNIDV_RANGE          
`define REQ_FLIT_STASHLPIDVALID_RANGE   `DSU_CHI_REQ_FLIT_STASHLPIDVALID_RANGE               
`define REQ_FLIT_STASHLPID_RANGE        `DSU_CHI_REQ_FLIT_STASHLPID_RANGE          
`define REQ_FLIT_RETURNTXNID_RANGE      `DSU_CHI_REQ_FLIT_RETURNTXNID_RANGE            
`define REQ_FLIT_OPCODE_RANGE           `DSU_CHI_REQ_FLIT_OPCODE_RANGE       
`define REQ_FLIT_SIZE_RANGE             `DSU_CHI_REQ_FLIT_SIZE_RANGE     
`define REQ_FLIT_ADDR_RANGE             `DSU_CHI_REQ_FLIT_ADDR_RANGE     
`define REQ_FLIT_NS_RANGE               `DSU_CHI_REQ_FLIT_NS_RANGE   
`define REQ_FLIT_LS_RANGE               `DSU_CHI_REQ_FLIT_LS_RANGE   
`define REQ_FLIT_ALLOWRETRY_RANGE       `DSU_CHI_REQ_FLIT_ALLOWRETRY_RANGE           
`define REQ_FLIT_ORDER_RANGE            `DSU_CHI_REQ_FLIT_ORDER_RANGE      
`define REQ_FLIT_PCRDTYPE_RANGE         `DSU_CHI_REQ_FLIT_PCRDTYPE_RANGE         
`define REQ_FLIT_MEMATTR_RANGE          `DSU_CHI_REQ_FLIT_MEMATTR_RANGE        
`define REQ_FLIT_MEMATTREWACK_RANGE     `DSU_CHI_REQ_FLIT_MEMATTREWACK_RANGE             
`define REQ_FLIT_MEMATTRCACHE_RANGE     `DSU_CHI_REQ_FLIT_MEMATTRCACHE_RANGE             
`define REQ_FLIT_MEMATTRALLHINT_RANGE   `DSU_CHI_REQ_FLIT_MEMATTRALLHINT_RANGE               
`define REQ_FLIT_MEMATTRDEVICE_RANGE    `DSU_CHI_REQ_FLIT_MEMATTRDEVICE_RANGE              
`define REQ_FLIT_SNPATTR_RANGE          `DSU_CHI_REQ_FLIT_SNPATTR_RANGE        
`define REQ_FLIT_LPID_RANGE             `DSU_CHI_REQ_FLIT_LPID_RANGE     
`define REQ_FLIT_EXCL_RANGE             `DSU_CHI_REQ_FLIT_EXCL_RANGE     
`define REQ_FLIT_EXPCOMPACK_RANGE       `DSU_CHI_REQ_FLIT_EXPCOMPACK_RANGE           
`define REQ_FLIT_TAGOP_RANGE            `DSU_CHI_REQ_FLIT_TAGOP_RANGE      
`define REQ_FLIT_TRACETAG_RANGE         `DSU_CHI_REQ_FLIT_TRACETAG_RANGE         
`define REQ_FLIT_MPAM_RANGE             `DSU_CHI_REQ_FLIT_MPAM_RANGE     
`define REQ_FLIT_RSVD_RANGE             `DSU_CHI_REQ_FLIT_RSVD_RANGE     
`define REQ_FLIT_SRCTYPE_RANGE          `DSU_CHI_REQ_FLIT_SRCTYPE_RANGE        
`define REQ_FLIT_LDID_RANGE             `DSU_CHI_REQ_FLIT_LDID_RANGE  

`define REQ_FLIT_QOS_WIDTH              `DSU_CHI_REQ_FLIT_QOS_WIDTH                  
`define REQ_FLIT_TGTID_WIDTH            `DSU_CHI_REQ_FLIT_TGTID_WIDTH                    
`define REQ_FLIT_SRCID_WIDTH            `DSU_CHI_REQ_FLIT_SRCID_WIDTH                    
`define REQ_FLIT_TXNID_WIDTH            `DSU_CHI_REQ_FLIT_TXNID_WIDTH                    
`define REQ_FLIT_RNID_WIDTH             `DSU_CHI_REQ_FLIT_RNID_WIDTH                   
`define REQ_FLIT_STASHNIDV_WIDTH        `DSU_CHI_REQ_FLIT_STASHNIDV_WIDTH                        
`define REQ_FLIT_RETURNTXNID_WIDTH      `DSU_CHI_REQ_FLIT_RETURNTXNID_WIDTH                          
`define REQ_FLIT_STASHLPID_WIDTH        `DSU_CHI_REQ_FLIT_STASHLPID_WIDTH                        
`define REQ_FLIT_STASHLPIDVALID_WIDTH   `DSU_CHI_REQ_FLIT_STASHLPIDVALID_WIDTH                             
`define REQ_FLIT_OPCODE_WIDTH           `DSU_CHI_REQ_FLIT_OPCODE_WIDTH                     
`define REQ_FLIT_SIZE_WIDTH             `DSU_CHI_REQ_FLIT_SIZE_WIDTH                   
`define REQ_FLIT_ADDR_WIDTH             `DSU_CHI_REQ_FLIT_ADDR_WIDTH                   
`define REQ_FLIT_NS_WIDTH               `DSU_CHI_REQ_FLIT_NS_WIDTH                 
`define REQ_FLIT_LS_WIDTH               `DSU_CHI_REQ_FLIT_LS_WIDTH                 
`define REQ_FLIT_ALLOWRETRY_WIDTH       `DSU_CHI_REQ_FLIT_ALLOWRETRY_WIDTH                         
`define REQ_FLIT_ORDER_WIDTH            `DSU_CHI_REQ_FLIT_ORDER_WIDTH                    
`define REQ_FLIT_PCRDTYPE_WIDTH         `DSU_CHI_REQ_FLIT_PCRDTYPE_WIDTH                       
`define REQ_FLIT_MEMATTR_WIDTH          `DSU_CHI_REQ_FLIT_MEMATTR_WIDTH                      
`define REQ_FLIT_MEMATTREWACK_WIDTH     `DSU_CHI_REQ_FLIT_MEMATTREWACK_WIDTH                           
`define REQ_FLIT_MEMATTRDEVICE_WIDTH    `DSU_CHI_REQ_FLIT_MEMATTRDEVICE_WIDTH                            
`define REQ_FLIT_MEMATTRCACHE_WIDTH     `DSU_CHI_REQ_FLIT_MEMATTRCACHE_WIDTH                           
`define REQ_FLIT_MEMATTRALLHINT_WIDTH   `DSU_CHI_REQ_FLIT_MEMATTRALLHINT_WIDTH                             
`define REQ_FLIT_SNPATTR_WIDTH          `DSU_CHI_REQ_FLIT_SNPATTR_WIDTH                      
`define REQ_FLIT_LPID_WIDTH             `DSU_CHI_REQ_FLIT_LPID_WIDTH                   
`define REQ_FLIT_EXCL_WIDTH             `DSU_CHI_REQ_FLIT_EXCL_WIDTH                   
`define REQ_FLIT_EXPCOMPACK_WIDTH       `DSU_CHI_REQ_FLIT_EXPCOMPACK_WIDTH                         
`define REQ_FLIT_TAGOP_WIDTH            `DSU_CHI_REQ_FLIT_TAGOP_WIDTH                    
`define REQ_FLIT_TRACETAG_WIDTH         `DSU_CHI_REQ_FLIT_TRACETAG_WIDTH                       
`define REQ_FLIT_MPAM_WIDTH             `DSU_CHI_REQ_FLIT_MPAM_WIDTH                   
`define REQ_FLIT_RSVD_WIDTH             `DSU_CHI_REQ_FLIT_RSVD_WIDTH                   
`define REQ_FLIT_SRCTYPE_WIDTH          `DSU_CHI_REQ_FLIT_SRCTYPE_WIDTH                      
`define REQ_FLIT_LDID_WIDTH             `DSU_CHI_REQ_FLIT_LDID_WIDTH                   

/*RSP FLIT*/
//CHI B
// `define RSP_FLIT_QOS_RANGE           `DSU_CHI_RSP_FLIT_QOS_RANGE
// `define RSP_FLIT_TGTID_RANGE         `DSU_CHI_RSP_FLIT_TGTID_RANGE
// `define RSP_FLIT_SRCID_RANGE         `DSU_CHI_RSP_FLIT_SRCID_RANGE
// `define RSP_FLIT_TXNID_RANGE         `DSU_CHI_RSP_FLIT_TXNID_RANGE
// `define RSP_FLIT_OPCODE_RANGE        `DSU_CHI_RSP_FLIT_OPCODE_RANGE
// `define RSP_FLIT_RESPERR_RANGE       `DSU_CHI_RSP_FLIT_RESPERR_RANGE
// `define RSP_FLIT_RESP_RANGE          `DSU_CHI_RSP_FLIT_RESP_RANGE
// `define RSP_FLIT_FWDSTATE_RANGE      `DSU_CHI_RSP_FLIT_FWDSTATE_RANGE
// `define RSP_FLIT_DBID_RANGE          `DSU_CHI_RSP_FLIT_DBID_RANGE
// `define RSP_FLIT_PCRDTYPE_RANGE      `DSU_CHI_RSP_FLIT_PCRDTYPE_RANGE
// `define RSP_FLIT_TRACETAG_RANGE      `DSU_CHI_RSP_FLIT_TRACETAG_RANGE
// `define RSP_FLIT_DEVEVENT_RANGE      `DSU_CHI_RSP_FLIT_DEVEVENT_RANGE

//CHI E
`define RSP_FLIT_QOS_RANGE              `DSU_CHI_RSP_FLIT_QOS_RANGE
`define RSP_FLIT_DEVICEID_RANGE         `DSU_CHI_RSP_FLIT_DEVICEID_RANGE     
`define RSP_FLIT_PORTID_RANGE           `DSU_CHI_RSP_FLIT_PORTID_RANGE   
`define RSP_FLIT_YID_RANGE              `DSU_CHI_RSP_FLIT_YID_RANGE
`define RSP_FLIT_XID_RANGE              `DSU_CHI_RSP_FLIT_XID_RANGE
`define RSP_FLIT_MESHID_RANGE           `DSU_CHI_RSP_FLIT_MESHID_RANGE   
`define RSP_FLIT_TGTID_RANGE            `DSU_CHI_RSP_FLIT_TGTID_RANGE  
`define RSP_FLIT_SRCID_RANGE            `DSU_CHI_RSP_FLIT_SRCID_RANGE  
`define RSP_FLIT_TXNID_RANGE            `DSU_CHI_RSP_FLIT_TXNID_RANGE  
`define RSP_FLIT_OPCODE_RANGE           `DSU_CHI_RSP_FLIT_OPCODE_RANGE   
`define RSP_FLIT_RESPERR_RANGE          `DSU_CHI_RSP_FLIT_RESPERR_RANGE    
`define RSP_FLIT_RESP_RANGE             `DSU_CHI_RSP_FLIT_RESP_RANGE 
`define RSP_FLIT_RESPSNP_RANGE          `DSU_CHI_RSP_FLIT_RESPSNP_RANGE    
`define RSP_FLIT_RESPPASSDIRTY_RANGE    `DSU_CHI_RSP_FLIT_RESPPASSDIRTY_RANGE          
`define RSP_FLIT_FWDSTATE_RANGE         `DSU_CHI_RSP_FLIT_FWDSTATE_RANGE     
`define RSP_FLIT_CBUSY_RANGE            `DSU_CHI_RSP_FLIT_CBUSY_RANGE  
`define RSP_FLIT_DBID_RANGE             `DSU_CHI_RSP_FLIT_DBID_RANGE 
`define RSP_FLIT_PCRDTYPE_RANGE         `DSU_CHI_RSP_FLIT_PCRDTYPE_RANGE     
`define RSP_FLIT_TAGOP_RANGE            `DSU_CHI_RSP_FLIT_TAGOP_RANGE  
`define RSP_FLIT_TRACETAG_RANGE         `DSU_CHI_RSP_FLIT_TRACETAG_RANGE     
`define RSP_FLIT_DEVEVENT_RANGE         `DSU_CHI_RSP_FLIT_DEVEVENT_RANGE 

`define RSP_FLIT_QOS_WIDTH             `DSU_CHI_RSP_FLIT_QOS_WIDTH  
`define RSP_FLIT_TGTID_WIDTH           `DSU_CHI_RSP_FLIT_TGTID_WIDTH    
`define RSP_FLIT_SRCID_WIDTH           `DSU_CHI_RSP_FLIT_SRCID_WIDTH    
`define RSP_FLIT_TXNID_WIDTH           `DSU_CHI_RSP_FLIT_TXNID_WIDTH    
`define RSP_FLIT_OPCODE_WIDTH          `DSU_CHI_RSP_FLIT_OPCODE_WIDTH     
`define RSP_FLIT_RESPERR_WIDTH         `DSU_CHI_RSP_FLIT_RESPERR_WIDTH      
`define RSP_FLIT_RESP_WIDTH            `DSU_CHI_RSP_FLIT_RESP_WIDTH   
`define RSP_FLIT_RESPSNP_WIDTH         `DSU_CHI_RSP_FLIT_RESPSNP_WIDTH      
`define RSP_FLIT_RESPPASSDIRTY_WIDTH   `DSU_CHI_RSP_FLIT_RESPPASSDIRTY_WIDTH            
`define RSP_FLIT_FWDSTATE_WIDTH        `DSU_CHI_RSP_FLIT_FWDSTATE_WIDTH       
`define RSP_FLIT_CBUSY_WIDTH           `DSU_CHI_RSP_FLIT_CBUSY_WIDTH    
`define RSP_FLIT_DBID_WIDTH            `DSU_CHI_RSP_FLIT_DBID_WIDTH   
`define RSP_FLIT_PCRDTYPE_WIDTH        `DSU_CHI_RSP_FLIT_PCRDTYPE_WIDTH       
`define RSP_FLIT_TAGOP_WIDTH           `DSU_CHI_RSP_FLIT_TAGOP_WIDTH    
`define RSP_FLIT_TRACETAG_WIDTH        `DSU_CHI_RSP_FLIT_TRACETAG_WIDTH       
`define RSP_FLIT_DEVEVENT_WIDTH        `DSU_CHI_RSP_FLIT_DEVEVENT_WIDTH  

/*DAT FLIT*/
//CHI B
// `define DAT_FLIT_QOS_RANGE           `DSU_CHI_DAT_FLIT_QOS_RANGE
// `define DAT_FLIT_TGTID_RANGE         `DSU_CHI_DAT_FLIT_TGTID_RANGE
// `define DAT_FLIT_SRCID_RANGE         `DSU_CHI_DAT_FLIT_SRCID_RANGE
// `define DAT_FLIT_TXNID_RANGE         `DSU_CHI_DAT_FLIT_TXNID_RANGE
// `define DAT_FLIT_HNID_RANGE          `DSU_CHI_DAT_FLIT_HNID_RANGE
// `define DAT_FLIT_OPCODE_RANGE        `DSU_CHI_DAT_FLIT_OPCODE_RANGE
// `define DAT_FLIT_RESPERR_RANGE       `DSU_CHI_DAT_FLIT_RESPERR_RANGE
// `define DAT_FLIT_RESP_RANGE          `DSU_CHI_DAT_FLIT_RESP_RANGE
// `define DAT_FLIT_FWDSTATE_RANGE      `DSU_CHI_DAT_FLIT_FWDSTATE_RANGE
// `define DAT_FLIT_DBID_RANGE          `DSU_CHI_DAT_FLIT_DBID_RANGE
// `define DAT_FLIT_CCID_RANGE          `DSU_CHI_DAT_FLIT_CCID_RANGE
// `define DAT_FLIT_DATAID_RANGE        `DSU_CHI_DAT_FLIT_DATAID_RANGE
// `define DAT_FLIT_TRACETAG_RANGE      `DSU_CHI_DAT_FLIT_TRACETAG_RANGE
// `define DAT_FLIT_RSVD_RANGE          `DSU_CHI_DAT_FLIT_RSVD_RANGE
// `define DAT_FLIT_BE_RANGE            `DSU_CHI_DAT_FLIT_BE_RANGE
// `define DAT_FLIT_DATA_RANGE          `DSU_CHI_DAT_FLIT_DATA_RANGE
// `define DAT_FLIT_POISON_RANGE        `DSU_CHI_DAT_FLIT_POISON_RANGE
// `define DAT_FLIT_CHUNKV_RANGE        `DSU_CHI_DAT_FLIT_CHUNKV_RANGE
// `define DAT_FLIT_DEVEVENT_RANGE      `DSU_CHI_DAT_FLIT_DEVEVENT_RANGE

//CHI E
`define DAT_FLIT_QOS_RANGE              `DSU_CHI_DAT_FLIT_QOS_RANGE   
`define DAT_FLIT_DEVICEID_RANGE         `DSU_CHI_DAT_FLIT_DEVICEID_RANGE        
`define DAT_FLIT_PORTID_RANGE           `DSU_CHI_DAT_FLIT_PORTID_RANGE      
`define DAT_FLIT_YID_RANGE              `DSU_CHI_DAT_FLIT_YID_RANGE   
`define DAT_FLIT_XID_RANGE              `DSU_CHI_DAT_FLIT_XID_RANGE   
`define DAT_FLIT_MESHID_RANGE           `DSU_CHI_DAT_FLIT_MESHID_RANGE      
`define DAT_FLIT_TGTID_RANGE            `DSU_CHI_DAT_FLIT_TGTID_RANGE     
`define DAT_FLIT_SRCID_RANGE            `DSU_CHI_DAT_FLIT_SRCID_RANGE     
`define DAT_FLIT_TXNID_RANGE            `DSU_CHI_DAT_FLIT_TXNID_RANGE     
`define DAT_FLIT_HNID_RANGE             `DSU_CHI_DAT_FLIT_HNID_RANGE    
`define DAT_FLIT_OPCODE_RANGE           `DSU_CHI_DAT_FLIT_OPCODE_RANGE      
`define DAT_FLIT_RESPERR_RANGE          `DSU_CHI_DAT_FLIT_RESPERR_RANGE       
`define DAT_FLIT_RESP_RANGE             `DSU_CHI_DAT_FLIT_RESP_RANGE    
`define DAT_FLIT_FWDSTATE_RANGE         `DSU_CHI_DAT_FLIT_FWDSTATE_RANGE        
`define DAT_FLIT_CBUSY_RANGE            `DSU_CHI_DAT_FLIT_CBUSY_RANGE     
`define DAT_FLIT_DBID_RANGE             `DSU_CHI_DAT_FLIT_DBID_RANGE    
`define DAT_FLIT_CCID_RANGE             `DSU_CHI_DAT_FLIT_CCID_RANGE    
`define DAT_FLIT_DATAID_RANGE           `DSU_CHI_DAT_FLIT_DATAID_RANGE      
`define DAT_FLIT_TAGOP_RANGE            `DSU_CHI_DAT_FLIT_TAGOP_RANGE     
`define DAT_FLIT_TAG_RANGE              `DSU_CHI_DAT_FLIT_TAG_RANGE   
`define DAT_FLIT_TU_RANGE               `DSU_CHI_DAT_FLIT_TU_RANGE  
`define DAT_FLIT_TRACETAG_RANGE         `DSU_CHI_DAT_FLIT_TRACETAG_RANGE        
`define DAT_FLIT_RSVD_RANGE             `DSU_CHI_DAT_FLIT_RSVD_RANGE    
`define DAT_FLIT_BE_RANGE               `DSU_CHI_DAT_FLIT_BE_RANGE  
`define DAT_FLIT_DATA_RANGE             `DSU_CHI_DAT_FLIT_DATA_RANGE    
`define DAT_FLIT_DATACHECK_RANGE        `DSU_CHI_DAT_FLIT_DATACHECK_RANGE         
`define DAT_FLIT_POISON_RANGE           `DSU_CHI_DAT_FLIT_POISON_RANGE      
`define DAT_FLIT_CHUNKV_RANGE           `DSU_CHI_DAT_FLIT_CHUNKV_RANGE      
`define DAT_FLIT_DEVEVENT_RANGE         `DSU_CHI_DAT_FLIT_DEVEVENT_RANGE   

`define DAT_FLIT_QOS_WIDTH              `DSU_CHI_DAT_FLIT_QOS_WIDTH     
`define DAT_FLIT_TGTID_WIDTH            `DSU_CHI_DAT_FLIT_TGTID_WIDTH       
`define DAT_FLIT_SRCID_WIDTH            `DSU_CHI_DAT_FLIT_SRCID_WIDTH       
`define DAT_FLIT_TXNID_WIDTH            `DSU_CHI_DAT_FLIT_TXNID_WIDTH       
`define DAT_FLIT_HNID_WIDTH             `DSU_CHI_DAT_FLIT_HNID_WIDTH      
`define DAT_FLIT_OPCODE_WIDTH           `DSU_CHI_DAT_FLIT_OPCODE_WIDTH        
`define DAT_FLIT_RESPERR_WIDTH          `DSU_CHI_DAT_FLIT_RESPERR_WIDTH         
`define DAT_FLIT_RESP_WIDTH             `DSU_CHI_DAT_FLIT_RESP_WIDTH      
`define DAT_FLIT_FWDSTATE_WIDTH         `DSU_CHI_DAT_FLIT_FWDSTATE_WIDTH          
`define DAT_FLIT_CBUSY_WIDTH            `DSU_CHI_DAT_FLIT_CBUSY_WIDTH       
`define DAT_FLIT_DBID_WIDTH             `DSU_CHI_DAT_FLIT_DBID_WIDTH      
`define DAT_FLIT_CCID_WIDTH             `DSU_CHI_DAT_FLIT_CCID_WIDTH      
`define DAT_FLIT_DATAID_WIDTH           `DSU_CHI_DAT_FLIT_DATAID_WIDTH        
`define DAT_FLIT_TAGOP_WIDTH            `DSU_CHI_DAT_FLIT_TAGOP_WIDTH       
`define DAT_FLIT_TAG_WIDTH              `DSU_CHI_DAT_FLIT_TAG_WIDTH     
`define DAT_FLIT_TU_WIDTH               `DSU_CHI_DAT_FLIT_TU_WIDTH    
`define DAT_FLIT_TRACETAG_WIDTH         `DSU_CHI_DAT_FLIT_TRACETAG_WIDTH          
`define DAT_FLIT_RSVD_WIDTH             `DSU_CHI_DAT_FLIT_RSVD_WIDTH      
`define DAT_FLIT_BE_WIDTH               `DSU_CHI_DAT_FLIT_BE_WIDTH    
`define DAT_FLIT_DATA_WIDTH             `DSU_CHI_DAT_FLIT_DATA_WIDTH      
`define DAT_FLIT_DATACHECK_WIDTH        `DSU_CHI_DAT_FLIT_DATACHECK_WIDTH           
`define DAT_FLIT_POISON_WIDTH           `DSU_CHI_DAT_FLIT_POISON_WIDTH        
`define DAT_FLIT_CHUNKV_WIDTH           `DSU_CHI_DAT_FLIT_CHUNKV_WIDTH        
`define DAT_FLIT_DEVEVENT_WIDTH         `DSU_CHI_DAT_FLIT_DEVEVENT_WIDTH          


/*SNP FLIT*/
//CHI B
// `define SNP_FLIT_QOS_RANGE           `DSU_CHI_SNP_FLIT_QOS_RANGE
// `define SNP_FLIT_SRCID_RANGE         `DSU_CHI_SNP_FLIT_SRCID_RANGE
// `define SNP_FLIT_TXNID_RANGE         `DSU_CHI_SNP_FLIT_TXNID_RANGE
// `define SNP_FLIT_FWDNID_RANGE        `DSU_CHI_SNP_FLIT_FWDNID_RANGE
// `define SNP_FLIT_FWDTXNID_RANGE      `DSU_CHI_SNP_FLIT_FWDTXNID_RANGE
// `define SNP_FLIT_OPCODE_RANGE        `DSU_CHI_SNP_FLIT_OPCODE_RANGE
// `define SNP_FLIT_ADDR_RANGE          `DSU_CHI_SNP_FLIT_ADDR_RANGE
// `define SNP_FLIT_NS_RANGE            `DSU_CHI_SNP_FLIT_NS_RANGE
// `define SNP_FLIT_DONOTGOTOSD_RANGE   `DSU_CHI_SNP_FLIT_DONOTGOTOSD_RANGE
// `define SNP_FLIT_RETTO_SRC_RANGE     `DSU_CHI_SNP_FLIT_RETTO_SRC_RANGE
// `define SNP_FLIT_TRACETAG_RANGE      `DSU_CHI_SNP_FLIT_TRACETAG_RANGE
// `define SNP_FLIT_LDID_RANGE          `DSU_CHI_SNP_FLIT_LDID_RANGE
// `define SNP_FLIT_TGTID_RANGE         `DSU_CHI_SNP_FLIT_TGTID_RANGE

//CHI E
`define SNP_FLIT_QOS_RANGE           `DSU_CHI_SNP_FLIT_QOS_RANGE   
`define SNP_FLIT_SRCID_RANGE         `DSU_CHI_SNP_FLIT_SRCID_RANGE     
`define SNP_FLIT_TXNID_RANGE         `DSU_CHI_SNP_FLIT_TXNID_RANGE     
`define SNP_FLIT_FWDNID_RANGE        `DSU_CHI_SNP_FLIT_FWDNID_RANGE      
`define SNP_FLIT_FWDTXNID_RANGE      `DSU_CHI_SNP_FLIT_FWDTXNID_RANGE        
`define SNP_FLIT_OPCODE_RANGE        `DSU_CHI_SNP_FLIT_OPCODE_RANGE      
`define SNP_FLIT_ADDR_RANGE          `DSU_CHI_SNP_FLIT_ADDR_RANGE    
`define SNP_FLIT_NS_RANGE            `DSU_CHI_SNP_FLIT_NS_RANGE  
`define SNP_FLIT_DONOTGOTOSD_RANGE   `DSU_CHI_SNP_FLIT_DONOTGOTOSD_RANGE           
`define SNP_FLIT_RETTO_SRC_RANGE     `DSU_CHI_SNP_FLIT_RETTO_SRC_RANGE         
`define SNP_FLIT_TRACETAG_RANGE      `DSU_CHI_SNP_FLIT_TRACETAG_RANGE        
`define SNP_FLIT_MPAM_RANGE          `DSU_CHI_SNP_FLIT_MPAM_RANGE    
`define SNP_FLIT_LDID_RANGE          `DSU_CHI_SNP_FLIT_LDID_RANGE    
`define SNP_FLIT_DEVICEID_RANGE      `DSU_CHI_SNP_FLIT_DEVICEID_RANGE        
`define SNP_FLIT_PORTID_RANGE        `DSU_CHI_SNP_FLIT_PORTID_RANGE      
`define SNP_FLIT_YID_RANGE           `DSU_CHI_SNP_FLIT_YID_RANGE   
`define SNP_FLIT_XID_RANGE           `DSU_CHI_SNP_FLIT_XID_RANGE   
`define SNP_FLIT_MESHID_RANGE        `DSU_CHI_SNP_FLIT_MESHID_RANGE      
`define SNP_FLIT_TGTID_RANGE         `DSU_CHI_SNP_FLIT_TGTID_RANGE 

`define SNP_FLIT_QOS_WIDTH           `DSU_CHI_SNP_FLIT_QOS_WIDTH 
`define SNP_FLIT_SRCID_WIDTH         `DSU_CHI_SNP_FLIT_SRCID_WIDTH   
`define SNP_FLIT_TXNID_WIDTH         `DSU_CHI_SNP_FLIT_TXNID_WIDTH   
`define SNP_FLIT_FWDNID_WIDTH        `DSU_CHI_SNP_FLIT_FWDNID_WIDTH    
`define SNP_FLIT_FWDTXNID_WIDTH      `DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH      
`define SNP_FLIT_OPCODE_WIDTH        `DSU_CHI_SNP_FLIT_OPCODE_WIDTH    
`define SNP_FLIT_ADDR_WIDTH          `DSU_CHI_SNP_FLIT_ADDR_WIDTH  
`define SNP_FLIT_NS_WIDTH            `DSU_CHI_SNP_FLIT_NS_WIDTH
`define SNP_FLIT_DONOTGOTOSD_WIDTH   `DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH         
`define SNP_FLIT_RETTO_SRC_WIDTH     `DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH       
`define SNP_FLIT_TRACETAG_WIDTH      `DSU_CHI_SNP_FLIT_TRACETAG_WIDTH      
`define SNP_FLIT_MPAM_WIDTH          `DSU_CHI_SNP_FLIT_MPAM_WIDTH  
`define SNP_FLIT_LDID_WIDTH          `DSU_CHI_SNP_FLIT_LDID_WIDTH  
`define SNP_FLIT_TGTID_WIDTH         `DSU_CHI_SNP_FLIT_TGTID_WIDTH   

/*DLB HEADER FLIT*/
`define DLB_FLIT_OPCODE_RANGE        `DSU_DLB_MESH_OPCODE_RANGE
`define DLB_FLIT_DEVICEID_RANGE      `DSU_DLB_MESH_DEVICEID_RANGE
`define DLB_FLIT_PORTID_RANGE        `DSU_DLB_MESH_PORTID_RANGE
`define DLB_FLIT_TODEV_RANGE         `DSU_DLB_MESH_TODEV_RANGE
`define DLB_FLIT_YID_RANGE           `DSU_DLB_MESH_YID_RANGE
`define DLB_FLIT_XID_RANGE           `DSU_DLB_MESH_XID_RANGE
`define DLB_FLIT_TGTID_RANGE         `DSU_DLB_MESH_TGTID_RANGE
`define DLB_FLIT_BRDCST_RANGE        `DSU_DLB_MESH_BRDCST_RANGE
`define DLB_FLIT_NEXT_RANGE          `DSU_DLB_NEXT_RANGE

//GLObAL SIGNAL
`define NOC_TLR_FLIT_WIDTH                    (`NOC_TLR_FLIT_RESET_WIDTH + `NOC_TLR_FLIT_DFTRSTDISABLE_WIDTH + `NOC_TLR_FLIT_SNAPSHOT_WIDTH)

`define NOC_TLR_FLIT_RESET_WIDTH              1
`define NOC_TLR_FLIT_DFTRSTDISABLE_WIDTH      1

`define NOC_TLR_FLIT_GLOBALSIG_WIDTH          (`NOC_TLR_FLIT_RESET_WIDTH + `NOC_TLR_FLIT_DFTRSTDISABLE_WIDTH)

`define NOC_TLR_FLIT_SNAPSHOT_VALID_WIDTH     1
`define NOC_TLR_FLIT_SNAPSHOT_FLIT_WIDTH      4

`define NOC_TLR_FLIT_SNAPSHOT_WIDTH           (`NOC_TLR_FLIT_SNAPSHOT_VALID_WIDTH + `NOC_TLR_FLIT_SNAPSHOT_FLIT_WIDTH)

`define NOC_TLR_FLIT_RESET_RIGHT              0
`define NOC_TLR_FLIT_RESET_LEFT               (`NOC_TLR_FLIT_RESET_RIGHT + `NOC_TLR_FLIT_RESET_WIDTH -1)
`define NOC_TLR_FLIT_DFTRSTDISABLE_RIGHT      (`NOC_TLR_FLIT_RESET_LEFT + 1)
`define NOC_TLR_FLIT_DFTRSTDISABLE_LEFT       (`NOC_TLR_FLIT_DFTRSTDISABLE_RIGHT + `NOC_TLR_FLIT_DFTRSTDISABLE_WIDTH -1)

`define NOC_TLR_FLIT_SNAPSHOT_VALID_RIGHT     (`NOC_TLR_FLIT_DFTRSTDISABLE_LEFT +1)
`define NOC_TLR_FLIT_SNAPSHOT_VALID_LEFT      (`NOC_TLR_FLIT_SNAPSHOT_VALID_RIGHT + `NOC_TLR_FLIT_SNAPSHOT_VALID_WIDTH-1)
`define NOC_TLR_FLIT_SNAPSHOT_FLIT_RIGHT      (`NOC_TLR_FLIT_SNAPSHOT_VALID_LEFT + 1)
`define NOC_TLR_FLIT_SNAPSHOT_FLIT_LEFT       (`NOC_TLR_FLIT_SNAPSHOT_FLIT_RIGHT + `NOC_TLR_FLIT_SNAPSHOT_FLIT_WIDTH-1)

`define NOC_TLR_FLIT_RESET_RANGE             `NOC_TLR_FLIT_RESET_LEFT  : `NOC_TLR_FLIT_RESET_RIGHT 
`define NOC_TLR_FLIT_DFTRSTDISABLE_RANGE     `NOC_TLR_FLIT_DFTRSTDISABLE_LEFT  : `NOC_TLR_FLIT_DFTRSTDISABLE_RIGHT 
`define NOC_TLR_FLIT_SNAPSHOT_VALID_RANGE    `NOC_TLR_FLIT_SNAPSHOT_VALID_LEFT : `NOC_TLR_FLIT_SNAPSHOT_VALID_RIGHT
`define NOC_TLR_FLIT_SNAPSHOT_FLIT_RANGE     `NOC_TLR_FLIT_SNAPSHOT_FLIT_LEFT  : `NOC_TLR_FLIT_SNAPSHOT_FLIT_RIGHT 

`define NOC_SNAPSHOT                         1

`define NOC_TLR_FLIT_INIT_VALUE              {5'b00000, 1'b0, 1'b0}

/*RNSAM*/
`define PA_RANGE                     `DSU_CHI_REQ_FLIT_ADDR_WIDTH-1 : 0
`define PA_WIDTH                     `DSU_CHI_REQ_FLIT_ADDR_WIDTH
`define NOC_NODEID_WIDTH             `DSU_NODEID_WIDTH

`define HNF_NID_W                    `DSU_NODEID_WIDTH

`define BASE_ADDR0                   `DSU_BASE_ADDR0
`define BASE_ADDR0_OFFSET            `DSU_BASE_ADDR0_OFFSET

`define BASE_ADDR1                   `DSU_BASE_ADDR1
`define BASE_ADDR1_OFFSET            `DSU_BASE_ADDR1_OFFSET

`define DEV_TYPE_RNFBESAM            `DSU_DEV_TYPE_RNFBESAM 
`define DEV_TYPE_SNF                 `DSU_DEV_TYPE_SNF     
`define DEV_TYPE_RNI                 `DSU_DEV_TYPE_RNI     
`define DEV_TYPE_OTHERS              `DSU_DEV_TYPE_OTHERS  

`define NONHASH_NODEID_WIDTH         16
`define NONHASH_NODE_VALID_RANGE     15:15
`define NONHASH_NODE_DEV_TYPE_RANGE  14:11
`define NONHASH_NODE_TGTID_RANGE     10:0

/*MDL*/
`define NOC_MDL_CHI_DEV0             0
`define NOC_MDL_CHI_DEV1             1
`define NOC_MDL_CHI_DEV2             2
`define NOC_MDL_CHI_DEV3             3

`define NOC_MDL_DLB_RUT              0
`define NOC_MDL_DLB_DEV0             1
`define NOC_MDL_DLB_DEV1             2
`define NOC_MDL_DLB_DEV2             3
`define NOC_MDL_DLB_DEV3             4

/*OTHER*/
`define NOC_LDID_WIDTH               `DSU_CHI_REQ_FLIT_LDID_WIDTH
`define NOC_DELAY                    0.1
`define NOC_LAT_DELAY                0
