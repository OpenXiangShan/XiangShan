//------------------------------------------------------------------------------
/*
    Copyright all by the Beijing Institute of Open Source CHIBip

    Filename    : dsu_chie_defines.sv
    File-history: 
       (1) Junyan Xie created on 2025/04/03 as the CHI-E-related macro definition file

  */

// TX Channel Handshake Signals
`define DSU_CHI_TX_LINKACTIVEREQ              1  // Placeholder value
`define DSU_CHI_TX_LINKACTIVEACK              1  // Placeholder value

// RX Channel Handshake Signals
`define DSU_CHI_RX_LINKACTIVEREQ              1  // Placeholder value
`define DSU_CHI_RX_LINKACTIVEACK              1  // Placeholder value

//NODEID
`define DSU_NODEID_WIDTH                       (0 + `DSU_MXP_DEVICEID_WIDTH_PARAM + `DSU_MXP_PORTID_WIDTH_PARAM + `DSU_MXP_YID_WIDTH_PARAM + `DSU_MXP_XID_WIDTH_PARAM + `DSU_MXP_MESHID_WIDTH_PARAM)
`define DSU_MXP_DEVICEID_WIDTH_PARAM           2
`define DSU_MXP_PORTID_WIDTH_PARAM             2
`define DSU_MXP_MESHID_WIDTH_PARAM             0
`define DSU_MXP_XID_WIDTH_PARAM                4
`define DSU_MXP_YID_WIDTH_PARAM                3

`define DSU_CHI_REQ_FLIT_QOS_WIDTH            4   //3:0
`define DSU_CHI_REQ_FLIT_TGTID_WIDTH          `DSU_NODEID_WIDTH //14:4
`define DSU_CHI_REQ_FLIT_SRCID_WIDTH          `DSU_NODEID_WIDTH //25:15   
`define DSU_CHI_REQ_FLIT_TXNID_WIDTH          12  //37:26
`define DSU_CHI_REQ_FLIT_RNID_WIDTH           `DSU_NODEID_WIDTH //48:38
`define DSU_CHI_REQ_FLIT_STASHNIDV_WIDTH      1   //49:49
`define DSU_CHI_REQ_FLIT_RETURNTXNID_WIDTH    12  //61:50
`define DSU_CHI_REQ_FLIT_STASHLPID_WIDTH      5   //54:50
`define DSU_CHI_REQ_FLIT_STASHLPIDVALID_WIDTH 1   //55:55
`define DSU_CHI_REQ_FLIT_OPCODE_WIDTH         7   //68:62
`define DSU_CHI_REQ_FLIT_SIZE_WIDTH           3   //71:69
`define DSU_CHI_REQ_FLIT_ADDR_WIDTH           48  //119:72
`define DSU_CHI_REQ_FLIT_NS_WIDTH             1   //120:120
`define DSU_CHI_REQ_FLIT_LS_WIDTH             1   //121:121
`define DSU_CHI_REQ_FLIT_ALLOWRETRY_WIDTH     1   //122:122
`define DSU_CHI_REQ_FLIT_ORDER_WIDTH          2   //124:123
`define DSU_CHI_REQ_FLIT_PCRDTYPE_WIDTH       4   //128:125
`define DSU_CHI_REQ_FLIT_MEMATTR_WIDTH        (`DSU_CHI_REQ_FLIT_MEMATTREWACK_WIDTH + `DSU_CHI_REQ_FLIT_MEMATTRDEVICE_WIDTH + `DSU_CHI_REQ_FLIT_MEMATTRCACHE_WIDTH + `DSU_CHI_REQ_FLIT_MEMATTRALLHINT_WIDTH)   //132:129
`define DSU_CHI_REQ_FLIT_MEMATTREWACK_WIDTH   1   //129:129
`define DSU_CHI_REQ_FLIT_MEMATTRDEVICE_WIDTH  1   //130:130
`define DSU_CHI_REQ_FLIT_MEMATTRCACHE_WIDTH   1   //131:131 
`define DSU_CHI_REQ_FLIT_MEMATTRALLHINT_WIDTH 1   //132:132
`define DSU_CHI_REQ_FLIT_SNPATTR_WIDTH        1   //133:133
`define DSU_CHI_REQ_FLIT_LPID_WIDTH           8   //141:134
`define DSU_CHI_REQ_FLIT_EXCL_WIDTH           1   //142:142
`define DSU_CHI_REQ_FLIT_EXPCOMPACK_WIDTH     1   //143:143
`define DSU_CHI_REQ_FLIT_TAGOP_WIDTH          2   //145:144
`define DSU_CHI_REQ_FLIT_TRACETAG_WIDTH       1   //146:146
`define DSU_CHI_REQ_FLIT_MPAM_WIDTH           11  //157:147
`define DSU_CHI_REQ_FLIT_RSVD_WIDTH           4   //161:158
`define DSU_CHI_REQ_FLIT_SRCTYPE_WIDTH        4   //165:162
`define DSU_CHI_REQ_FLIT_LDID_WIDTH           6   //171:166


`define DSU_CHI_RSP_FLIT_QOS_WIDTH            4   //3:0
`define DSU_CHI_RSP_FLIT_TGTID_WIDTH          `DSU_NODEID_WIDTH   //14:4
`define DSU_CHI_RSP_FLIT_SRCID_WIDTH          `DSU_NODEID_WIDTH   //25:15   
`define DSU_CHI_RSP_FLIT_TXNID_WIDTH          12  //37:26
`define DSU_CHI_RSP_FLIT_OPCODE_WIDTH         5   //42:38 
`define DSU_CHI_RSP_FLIT_RESPERR_WIDTH        2   //44:43
`define DSU_CHI_RSP_FLIT_RESP_WIDTH           (`DSU_CHI_RSP_FLIT_RESPSNP_WIDTH + `DSU_CHI_RSP_FLIT_RESPPASSDIRTY_WIDTH)   //47:45
`define DSU_CHI_RSP_FLIT_RESPSNP_WIDTH        2   //46:45
`define DSU_CHI_RSP_FLIT_RESPPASSDIRTY_WIDTH  1   //47:47
`define DSU_CHI_RSP_FLIT_FWDSTATE_WIDTH       3   //50:48
`define DSU_CHI_RSP_FLIT_CBUSY_WIDTH          3   //53:51
`define DSU_CHI_RSP_FLIT_DBID_WIDTH           12  //65:54
`define DSU_CHI_RSP_FLIT_PCRDTYPE_WIDTH       4   //69:66
`define DSU_CHI_RSP_FLIT_TAGOP_WIDTH          2   //71:70
`define DSU_CHI_RSP_FLIT_TRACETAG_WIDTH       1   //72:72
`define DSU_CHI_RSP_FLIT_DEVEVENT_WIDTH       2   //74:73


`define DSU_CHI_DAT_FLIT_QOS_WIDTH            4   //3:0   
`define DSU_CHI_DAT_FLIT_TGTID_WIDTH          `DSU_NODEID_WIDTH   //14:4
`define DSU_CHI_DAT_FLIT_SRCID_WIDTH          `DSU_NODEID_WIDTH   //25:15   
`define DSU_CHI_DAT_FLIT_TXNID_WIDTH          12  //37:26   
`define DSU_CHI_DAT_FLIT_HNID_WIDTH           `DSU_NODEID_WIDTH   //48:38 
`define DSU_CHI_DAT_FLIT_OPCODE_WIDTH         4   //52:49
`define DSU_CHI_DAT_FLIT_RESPERR_WIDTH        2   //54:53
`define DSU_CHI_DAT_FLIT_RESP_WIDTH           `DSU_CHI_RSP_FLIT_RESP_WIDTH  //57:55
`define DSU_CHI_DAT_FLIT_FWDSTATE_WIDTH       4   //61:58
`define DSU_CHI_DAT_FLIT_CBUSY_WIDTH          3   //64:62
`define DSU_CHI_DAT_FLIT_DBID_WIDTH           12  //76:65
`define DSU_CHI_DAT_FLIT_CCID_WIDTH           2   //78:77
`define DSU_CHI_DAT_FLIT_DATAID_WIDTH         2   //80:79
`define DSU_CHI_DAT_FLIT_TAGOP_WIDTH          2   //82:81
`define DSU_CHI_DAT_FLIT_TAG_WIDTH            8   //90:83
`define DSU_CHI_DAT_FLIT_TU_WIDTH             2   //92:91
`define DSU_CHI_DAT_FLIT_TRACETAG_WIDTH       1   //93:93
`define DSU_CHI_DAT_FLIT_RSVD_WIDTH           4   //97:94
`define DSU_CHI_DAT_FLIT_BE_WIDTH             32  //129:98
`define DSU_CHI_DAT_FLIT_DATA_WIDTH           256 //385:130
`define DSU_CHI_DAT_FLIT_DATACHECK_WIDTH      32  //417:386
`define DSU_CHI_DAT_FLIT_POISON_WIDTH         4   //421:418
`define DSU_CHI_DAT_FLIT_CHUNKV_WIDTH         2   //423:422
`define DSU_CHI_DAT_FLIT_DEVEVENT_WIDTH       2   //425:424


`define DSU_CHI_SNP_FLIT_QOS_WIDTH            4   //3:0
`define DSU_CHI_SNP_FLIT_SRCID_WIDTH          `DSU_NODEID_WIDTH   //14:4
`define DSU_CHI_SNP_FLIT_TXNID_WIDTH          12  //26:15
`define DSU_CHI_SNP_FLIT_FWDNID_WIDTH         `DSU_NODEID_WIDTH   //37:27   
`define DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH       12  //49:38
`define DSU_CHI_SNP_FLIT_OPCODE_WIDTH         5   //54:50
`define DSU_CHI_SNP_FLIT_ADDR_WIDTH           45  //99:55
`define DSU_CHI_SNP_FLIT_NS_WIDTH             1   //100:100
`define DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH    1   //101:101
`define DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH      1   //102:102
`define DSU_CHI_SNP_FLIT_TRACETAG_WIDTH       1   //103:103
`define DSU_CHI_SNP_FLIT_MPAM_WIDTH           11  //114:104
`define DSU_CHI_SNP_FLIT_LDID_WIDTH           6   //120:115
`define DSU_CHI_SNP_FLIT_TGTID_WIDTH          `DSU_NODEID_WIDTH //131:121


`define DSU_CHI_REQ_FLIT_WIDTH \
    (`DSU_CHI_REQ_FLIT_QOS_WIDTH + `DSU_CHI_REQ_FLIT_TGTID_WIDTH + `DSU_CHI_REQ_FLIT_SRCID_WIDTH + \
     `DSU_CHI_REQ_FLIT_TXNID_WIDTH + `DSU_CHI_REQ_FLIT_RNID_WIDTH + `DSU_CHI_REQ_FLIT_STASHNIDV_WIDTH + \
     `DSU_CHI_REQ_FLIT_RETURNTXNID_WIDTH + `DSU_CHI_REQ_FLIT_OPCODE_WIDTH + `DSU_CHI_REQ_FLIT_SIZE_WIDTH + \
     `DSU_CHI_REQ_FLIT_ADDR_WIDTH + `DSU_CHI_REQ_FLIT_NS_WIDTH + `DSU_CHI_REQ_FLIT_LS_WIDTH + \
     `DSU_CHI_REQ_FLIT_ALLOWRETRY_WIDTH + `DSU_CHI_REQ_FLIT_ORDER_WIDTH + `DSU_CHI_REQ_FLIT_PCRDTYPE_WIDTH + \
     `DSU_CHI_REQ_FLIT_MEMATTR_WIDTH + `DSU_CHI_REQ_FLIT_SNPATTR_WIDTH + `DSU_CHI_REQ_FLIT_LPID_WIDTH + \
     `DSU_CHI_REQ_FLIT_EXCL_WIDTH + `DSU_CHI_REQ_FLIT_EXPCOMPACK_WIDTH + `DSU_CHI_REQ_FLIT_TAGOP_WIDTH + \
     `DSU_CHI_REQ_FLIT_TRACETAG_WIDTH + `DSU_CHI_REQ_FLIT_MPAM_WIDTH + \
     `DSU_CHI_REQ_FLIT_RSVD_WIDTH + `DSU_CHI_REQ_FLIT_SRCTYPE_WIDTH + `DSU_CHI_REQ_FLIT_LDID_WIDTH)              

`define DSU_CHI_REQ_FLIT_RANGE                 (`DSU_CHI_REQ_FLIT_WIDTH-1) : 0         

`define DSU_CHI_RSP_FLIT_WIDTH \
    (`DSU_CHI_RSP_FLIT_QOS_WIDTH + `DSU_CHI_RSP_FLIT_TGTID_WIDTH + `DSU_CHI_RSP_FLIT_SRCID_WIDTH + \
     `DSU_CHI_RSP_FLIT_TXNID_WIDTH + `DSU_CHI_RSP_FLIT_OPCODE_WIDTH + `DSU_CHI_RSP_FLIT_RESPERR_WIDTH + \
     `DSU_CHI_RSP_FLIT_RESP_WIDTH + `DSU_CHI_RSP_FLIT_FWDSTATE_WIDTH + `DSU_CHI_RSP_FLIT_CBUSY_WIDTH + \
     `DSU_CHI_RSP_FLIT_DBID_WIDTH + `DSU_CHI_RSP_FLIT_PCRDTYPE_WIDTH + `DSU_CHI_RSP_FLIT_TAGOP_WIDTH + \
     `DSU_CHI_RSP_FLIT_TRACETAG_WIDTH + `DSU_CHI_RSP_FLIT_DEVEVENT_WIDTH)

`define DSU_CHI_RSP_FLIT_RANGE                 (`DSU_CHI_RSP_FLIT_WIDTH-1) : 0   

`define DSU_CHI_DAT_FLIT_WIDTH \
    (`DSU_CHI_DAT_FLIT_QOS_WIDTH + `DSU_CHI_DAT_FLIT_TGTID_WIDTH + `DSU_CHI_DAT_FLIT_SRCID_WIDTH + \
     `DSU_CHI_DAT_FLIT_TXNID_WIDTH + `DSU_CHI_DAT_FLIT_HNID_WIDTH + `DSU_CHI_DAT_FLIT_OPCODE_WIDTH + \
     `DSU_CHI_DAT_FLIT_RESPERR_WIDTH + `DSU_CHI_DAT_FLIT_RESP_WIDTH + `DSU_CHI_DAT_FLIT_FWDSTATE_WIDTH + \
     `DSU_CHI_DAT_FLIT_CBUSY_WIDTH + `DSU_CHI_DAT_FLIT_DBID_WIDTH + `DSU_CHI_DAT_FLIT_CCID_WIDTH + \
     `DSU_CHI_DAT_FLIT_DATAID_WIDTH + `DSU_CHI_DAT_FLIT_TAGOP_WIDTH + `DSU_CHI_DAT_FLIT_TAG_WIDTH + `DSU_CHI_DAT_FLIT_TU_WIDTH + \
     `DSU_CHI_DAT_FLIT_TRACETAG_WIDTH + `DSU_CHI_DAT_FLIT_RSVD_WIDTH + `DSU_CHI_DAT_FLIT_BE_WIDTH + \
     `DSU_CHI_DAT_FLIT_DATA_WIDTH + `DSU_CHI_DAT_FLIT_DATACHECK_WIDTH + `DSU_CHI_DAT_FLIT_POISON_WIDTH + \
     `DSU_CHI_DAT_FLIT_CHUNKV_WIDTH + `DSU_CHI_DAT_FLIT_DEVEVENT_WIDTH)

`define DSU_CHI_DAT_FLIT_RANGE                 (`DSU_CHI_DAT_FLIT_WIDTH-1) : 0   

`define DSU_CHI_SNP_FLIT_WIDTH \
    (`DSU_CHI_SNP_FLIT_QOS_WIDTH + `DSU_CHI_SNP_FLIT_SRCID_WIDTH + `DSU_CHI_SNP_FLIT_TXNID_WIDTH + \
     `DSU_CHI_SNP_FLIT_FWDNID_WIDTH + `DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH + `DSU_CHI_SNP_FLIT_OPCODE_WIDTH + \
     `DSU_CHI_SNP_FLIT_ADDR_WIDTH + `DSU_CHI_SNP_FLIT_NS_WIDTH + `DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH + \
     `DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH + `DSU_CHI_SNP_FLIT_TRACETAG_WIDTH + `DSU_CHI_SNP_FLIT_MPAM_WIDTH + \
     `DSU_CHI_SNP_FLIT_LDID_WIDTH + `DSU_CHI_SNP_FLIT_TGTID_WIDTH)

`define DSU_CHI_SNP_FLIT_RANGE                 (`DSU_CHI_SNP_FLIT_WIDTH-1) : 0   

`define DSU_CHI_SNP_FLIT_NO_TGTID_WIDTH \
    (`DSU_CHI_SNP_FLIT_QOS_WIDTH + `DSU_CHI_SNP_FLIT_SRCID_WIDTH + `DSU_CHI_SNP_FLIT_TXNID_WIDTH + \
     `DSU_CHI_SNP_FLIT_FWDNID_WIDTH + `DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH + `DSU_CHI_SNP_FLIT_OPCODE_WIDTH + \
     `DSU_CHI_SNP_FLIT_ADDR_WIDTH + `DSU_CHI_SNP_FLIT_NS_WIDTH + `DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH + \
     `DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH + `DSU_CHI_SNP_FLIT_TRACETAG_WIDTH + `DSU_CHI_SNP_FLIT_MPAM_WIDTH + \
     `DSU_CHI_SNP_FLIT_LDID_WIDTH)

`define DSU_CHI_SNP_FLIT_NO_TGTID_RANGE        (`DSU_CHI_SNP_FLIT_NO_TGTID_WIDTH-1) : 0

`define DSU_CHI_RNFBESAM_REQ_FLIT_WIDTH \
    (`DSU_CHI_REQ_FLIT_QOS_WIDTH + `DSU_CHI_REQ_FLIT_TGTID_WIDTH + `DSU_CHI_REQ_FLIT_SRCID_WIDTH + \
     `DSU_CHI_REQ_FLIT_TXNID_WIDTH + `DSU_CHI_REQ_FLIT_RNID_WIDTH + `DSU_CHI_REQ_FLIT_STASHNIDV_WIDTH + \
     `DSU_CHI_REQ_FLIT_RETURNTXNID_WIDTH + `DSU_CHI_REQ_FLIT_OPCODE_WIDTH + `DSU_CHI_REQ_FLIT_SIZE_WIDTH + \
     `DSU_CHI_REQ_FLIT_ADDR_WIDTH + `DSU_CHI_REQ_FLIT_NS_WIDTH + `DSU_CHI_REQ_FLIT_LS_WIDTH + \
     `DSU_CHI_REQ_FLIT_ALLOWRETRY_WIDTH + `DSU_CHI_REQ_FLIT_ORDER_WIDTH + `DSU_CHI_REQ_FLIT_PCRDTYPE_WIDTH + \
     `DSU_CHI_REQ_FLIT_MEMATTR_WIDTH + `DSU_CHI_REQ_FLIT_SNPATTR_WIDTH + `DSU_CHI_REQ_FLIT_LPID_WIDTH + \
     `DSU_CHI_REQ_FLIT_EXCL_WIDTH + `DSU_CHI_REQ_FLIT_EXPCOMPACK_WIDTH + `DSU_CHI_REQ_FLIT_TAGOP_WIDTH + \
     `DSU_CHI_REQ_FLIT_TRACETAG_WIDTH + `DSU_CHI_REQ_FLIT_MPAM_WIDTH + \
     `DSU_CHI_REQ_FLIT_RSVD_WIDTH)


`define DSU_CHI_RNFBESAM_RSP_FLIT_WIDTH \
    (`DSU_CHI_RSP_FLIT_QOS_WIDTH + `DSU_CHI_RSP_FLIT_TGTID_WIDTH + `DSU_CHI_RSP_FLIT_SRCID_WIDTH + \
     `DSU_CHI_RSP_FLIT_TXNID_WIDTH + `DSU_CHI_RSP_FLIT_OPCODE_WIDTH + `DSU_CHI_RSP_FLIT_RESPERR_WIDTH + \
     `DSU_CHI_RSP_FLIT_RESP_WIDTH + `DSU_CHI_RSP_FLIT_FWDSTATE_WIDTH + `DSU_CHI_RSP_FLIT_CBUSY_WIDTH + \
     `DSU_CHI_RSP_FLIT_DBID_WIDTH + `DSU_CHI_RSP_FLIT_PCRDTYPE_WIDTH + `DSU_CHI_RSP_FLIT_TAGOP_WIDTH + \
     `DSU_CHI_RSP_FLIT_TRACETAG_WIDTH)


`define DSU_CHI_RNFBESAM_SNP_FLIT_WIDTH \
    (`DSU_CHI_SNP_FLIT_QOS_WIDTH + `DSU_CHI_SNP_FLIT_SRCID_WIDTH + `DSU_CHI_SNP_FLIT_TXNID_WIDTH + \
     `DSU_CHI_SNP_FLIT_FWDNID_WIDTH + `DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH + `DSU_CHI_SNP_FLIT_OPCODE_WIDTH + \
     `DSU_CHI_SNP_FLIT_ADDR_WIDTH + `DSU_CHI_SNP_FLIT_NS_WIDTH + `DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH + \
     `DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH + `DSU_CHI_SNP_FLIT_TRACETAG_WIDTH + `DSU_CHI_SNP_FLIT_MPAM_WIDTH)


`define DSU_CHI_RNFBESAM_DAT_FLIT_WIDTH \
    (`DSU_CHI_DAT_FLIT_QOS_WIDTH + `DSU_CHI_DAT_FLIT_TGTID_WIDTH + `DSU_CHI_DAT_FLIT_SRCID_WIDTH + \
     `DSU_CHI_DAT_FLIT_TXNID_WIDTH + `DSU_CHI_DAT_FLIT_HNID_WIDTH + `DSU_CHI_DAT_FLIT_OPCODE_WIDTH + \
     `DSU_CHI_DAT_FLIT_RESPERR_WIDTH + `DSU_CHI_DAT_FLIT_RESP_WIDTH + `DSU_CHI_DAT_FLIT_FWDSTATE_WIDTH + \
     `DSU_CHI_DAT_FLIT_CBUSY_WIDTH + `DSU_CHI_DAT_FLIT_DBID_WIDTH + `DSU_CHI_DAT_FLIT_CCID_WIDTH + \
     `DSU_CHI_DAT_FLIT_DATAID_WIDTH + `DSU_CHI_DAT_FLIT_TAGOP_WIDTH + `DSU_CHI_DAT_FLIT_TAG_WIDTH + `DSU_CHI_DAT_FLIT_TU_WIDTH + \
     `DSU_CHI_DAT_FLIT_TRACETAG_WIDTH + `DSU_CHI_DAT_FLIT_RSVD_WIDTH + `DSU_CHI_DAT_FLIT_BE_WIDTH + \
     `DSU_CHI_DAT_FLIT_DATA_WIDTH + `DSU_CHI_DAT_FLIT_DATACHECK_WIDTH + `DSU_CHI_DAT_FLIT_POISON_WIDTH)


// Define the range parameterp
// QOS
`define DSU_CHI_REQ_FLIT_QOS_RIGHT    0
`define DSU_CHI_REQ_FLIT_QOS_LEFT     (`DSU_CHI_REQ_FLIT_QOS_RIGHT + `DSU_CHI_REQ_FLIT_QOS_WIDTH - 1)

// TGTID
`define DSU_CHI_REQ_FLIT_TGTID_RIGHT      (`DSU_CHI_REQ_FLIT_QOS_LEFT + 1)
`define DSU_CHI_REQ_FLIT_TGTID_LEFT       (`DSU_CHI_REQ_FLIT_TGTID_RIGHT + `DSU_CHI_REQ_FLIT_TGTID_WIDTH - 1)
`define DSU_CHI_REQ_FLIT_DEVICEID_RIGHT   (`DSU_CHI_REQ_FLIT_QOS_LEFT + 1)
`define DSU_CHI_REQ_FLIT_DEVICEID_LEFT    (`DSU_CHI_REQ_FLIT_DEVICEID_RIGHT + `DSU_MXP_DEVICEID_WIDTH_PARAM - 1)
`define DSU_CHI_REQ_FLIT_PORTID_RIGHT     (`DSU_CHI_REQ_FLIT_DEVICEID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_PORTID_LEFT      (`DSU_CHI_REQ_FLIT_PORTID_RIGHT + `DSU_MXP_PORTID_WIDTH_PARAM - 1)
`define DSU_CHI_REQ_FLIT_YID_RIGHT        (`DSU_CHI_REQ_FLIT_PORTID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_YID_LEFT         (`DSU_CHI_REQ_FLIT_YID_RIGHT + `DSU_MXP_YID_WIDTH_PARAM - 1)
`define DSU_CHI_REQ_FLIT_XID_RIGHT        (`DSU_CHI_REQ_FLIT_YID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_XID_LEFT         (`DSU_CHI_REQ_FLIT_XID_RIGHT + `DSU_MXP_XID_WIDTH_PARAM - 1)
`define DSU_CHI_REQ_FLIT_MESHID_RIGHT     (`DSU_CHI_REQ_FLIT_XID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MESHID_LEFT      (`DSU_CHI_REQ_FLIT_MESHID_RIGHT + `DSU_MXP_MESHID_WIDTH_PARAM - 1)

// SRCID
`define DSU_CHI_REQ_FLIT_SRCID_RIGHT  (`DSU_CHI_REQ_FLIT_TGTID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_SRCID_LEFT   (`DSU_CHI_REQ_FLIT_SRCID_RIGHT + `DSU_CHI_REQ_FLIT_SRCID_WIDTH - 1)

// TXNID
`define DSU_CHI_REQ_FLIT_TXNID_RIGHT  (`DSU_CHI_REQ_FLIT_SRCID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_TXNID_LEFT   (`DSU_CHI_REQ_FLIT_TXNID_RIGHT + `DSU_CHI_REQ_FLIT_TXNID_WIDTH - 1)

// RNID
`define DSU_CHI_REQ_FLIT_RNID_RIGHT   (`DSU_CHI_REQ_FLIT_TXNID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_RNID_LEFT    (`DSU_CHI_REQ_FLIT_RNID_RIGHT + `DSU_CHI_REQ_FLIT_RNID_WIDTH - 1)

// STASHNIDV
`define DSU_CHI_REQ_FLIT_STASHNIDV_RIGHT   (`DSU_CHI_REQ_FLIT_RNID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_STASHNIDV_LEFT    (`DSU_CHI_REQ_FLIT_STASHNIDV_RIGHT + `DSU_CHI_REQ_FLIT_STASHNIDV_WIDTH - 1)

// RETURNTXNID
`define DSU_CHI_REQ_FLIT_RETURNTXNID_RIGHT (`DSU_CHI_REQ_FLIT_STASHNIDV_LEFT + 1)
`define DSU_CHI_REQ_FLIT_RETURNTXNID_LEFT  (`DSU_CHI_REQ_FLIT_RETURNTXNID_RIGHT + `DSU_CHI_REQ_FLIT_RETURNTXNID_WIDTH - 1)

`define DSU_CHI_REQ_FLIT_STASHLPID_RIGHT   (`DSU_CHI_REQ_FLIT_STASHNIDV_LEFT + 1)
`define DSU_CHI_REQ_FLIT_STASHLPID_LEFT    (`DSU_CHI_REQ_FLIT_STASHLPID_RIGHT + `DSU_CHI_REQ_FLIT_STASHLPID_WIDTH - 1)   //addition

`define DSU_CHI_REQ_FLIT_STASHLPIDVALID_RIGHT (`DSU_CHI_REQ_FLIT_STASHLPID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_STASHLPIDVALID_LEFT  (`DSU_CHI_REQ_FLIT_STASHLPIDVALID_RIGHT + `DSU_CHI_REQ_FLIT_STASHLPIDVALID_WIDTH - 1) //addition


// OPCODE
`define DSU_CHI_REQ_FLIT_OPCODE_RIGHT  (`DSU_CHI_REQ_FLIT_RETURNTXNID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_OPCODE_LEFT   (`DSU_CHI_REQ_FLIT_OPCODE_RIGHT + `DSU_CHI_REQ_FLIT_OPCODE_WIDTH - 1)

// SIZE
`define DSU_CHI_REQ_FLIT_SIZE_RIGHT    (`DSU_CHI_REQ_FLIT_OPCODE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_SIZE_LEFT     (`DSU_CHI_REQ_FLIT_SIZE_RIGHT + `DSU_CHI_REQ_FLIT_SIZE_WIDTH - 1)

// ADDR
`define DSU_CHI_REQ_FLIT_ADDR_RIGHT    (`DSU_CHI_REQ_FLIT_SIZE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_ADDR_LEFT     (`DSU_CHI_REQ_FLIT_ADDR_RIGHT + `DSU_CHI_REQ_FLIT_ADDR_WIDTH - 1)

// NS
`define DSU_CHI_REQ_FLIT_NS_RIGHT      (`DSU_CHI_REQ_FLIT_ADDR_LEFT + 1)
`define DSU_CHI_REQ_FLIT_NS_LEFT       (`DSU_CHI_REQ_FLIT_NS_RIGHT + `DSU_CHI_REQ_FLIT_NS_WIDTH - 1)

// LS
`define DSU_CHI_REQ_FLIT_LS_RIGHT      (`DSU_CHI_REQ_FLIT_NS_LEFT + 1)
`define DSU_CHI_REQ_FLIT_LS_LEFT       (`DSU_CHI_REQ_FLIT_LS_RIGHT + `DSU_CHI_REQ_FLIT_LS_WIDTH - 1)

// ALLOWRETRY
`define DSU_CHI_REQ_FLIT_ALLOWRETRY_RIGHT  (`DSU_CHI_REQ_FLIT_LS_LEFT + 1)
`define DSU_CHI_REQ_FLIT_ALLOWRETRY_LEFT   (`DSU_CHI_REQ_FLIT_ALLOWRETRY_RIGHT + `DSU_CHI_REQ_FLIT_ALLOWRETRY_WIDTH - 1)

// ORDER
`define DSU_CHI_REQ_FLIT_ORDER_RIGHT   (`DSU_CHI_REQ_FLIT_ALLOWRETRY_LEFT + 1)
`define DSU_CHI_REQ_FLIT_ORDER_LEFT    (`DSU_CHI_REQ_FLIT_ORDER_RIGHT + `DSU_CHI_REQ_FLIT_ORDER_WIDTH - 1)

// PCRDTYPE
`define DSU_CHI_REQ_FLIT_PCRDTYPE_RIGHT    (`DSU_CHI_REQ_FLIT_ORDER_LEFT + 1)
`define DSU_CHI_REQ_FLIT_PCRDTYPE_LEFT     (`DSU_CHI_REQ_FLIT_PCRDTYPE_RIGHT + `DSU_CHI_REQ_FLIT_PCRDTYPE_WIDTH - 1)

// MEMATTR
`define DSU_CHI_REQ_FLIT_MEMATTR_RIGHT     (`DSU_CHI_REQ_FLIT_PCRDTYPE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MEMATTR_LEFT      (`DSU_CHI_REQ_FLIT_MEMATTR_RIGHT + `DSU_CHI_REQ_FLIT_MEMATTR_WIDTH - 1)

`define DSU_CHI_REQ_FLIT_MEMATTREWACK_RIGHT     (`DSU_CHI_REQ_FLIT_PCRDTYPE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MEMATTREWACK_LEFT      (`DSU_CHI_REQ_FLIT_MEMATTREWACK_RIGHT + `DSU_CHI_REQ_FLIT_MEMATTREWACK_WIDTH - 1)   

`define DSU_CHI_REQ_FLIT_MEMATTRDEVICE_RIGHT     (`DSU_CHI_REQ_FLIT_MEMATTREWACK_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MEMATTRDEVICE_LEFT      (`DSU_CHI_REQ_FLIT_MEMATTRDEVICE_RIGHT + `DSU_CHI_REQ_FLIT_MEMATTRDEVICE_WIDTH - 1)  

`define DSU_CHI_REQ_FLIT_MEMATTRCACHE_RIGHT     (`DSU_CHI_REQ_FLIT_MEMATTRDEVICE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MEMATTRCACHE_LEFT      (`DSU_CHI_REQ_FLIT_MEMATTRCACHE_RIGHT + `DSU_CHI_REQ_FLIT_MEMATTRCACHE_WIDTH - 1)  

`define DSU_CHI_REQ_FLIT_MEMATTRALLHINT_RIGHT     (`DSU_CHI_REQ_FLIT_MEMATTRCACHE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MEMATTRALLHINT_LEFT      (`DSU_CHI_REQ_FLIT_MEMATTRALLHINT_RIGHT + `DSU_CHI_REQ_FLIT_MEMATTRALLHINT_WIDTH - 1)  

// SNPATTR
`define DSU_CHI_REQ_FLIT_SNPATTR_RIGHT     (`DSU_CHI_REQ_FLIT_MEMATTR_LEFT + 1)
`define DSU_CHI_REQ_FLIT_SNPATTR_LEFT      (`DSU_CHI_REQ_FLIT_SNPATTR_RIGHT + `DSU_CHI_REQ_FLIT_SNPATTR_WIDTH - 1)

// LPID
`define DSU_CHI_REQ_FLIT_LPID_RIGHT        (`DSU_CHI_REQ_FLIT_SNPATTR_LEFT + 1)
`define DSU_CHI_REQ_FLIT_LPID_LEFT         (`DSU_CHI_REQ_FLIT_LPID_RIGHT + `DSU_CHI_REQ_FLIT_LPID_WIDTH - 1)

// EXCL
`define DSU_CHI_REQ_FLIT_EXCL_RIGHT        (`DSU_CHI_REQ_FLIT_LPID_LEFT + 1)
`define DSU_CHI_REQ_FLIT_EXCL_LEFT         (`DSU_CHI_REQ_FLIT_EXCL_RIGHT + `DSU_CHI_REQ_FLIT_EXCL_WIDTH - 1)

// EXPCOMPACK
`define DSU_CHI_REQ_FLIT_EXPCOMPACK_RIGHT  (`DSU_CHI_REQ_FLIT_EXCL_LEFT + 1)
`define DSU_CHI_REQ_FLIT_EXPCOMPACK_LEFT   (`DSU_CHI_REQ_FLIT_EXPCOMPACK_RIGHT + `DSU_CHI_REQ_FLIT_EXPCOMPACK_WIDTH - 1)

//TAGOP
`define DSU_CHI_REQ_FLIT_TAGOP_RIGHT       (`DSU_CHI_REQ_FLIT_EXPCOMPACK_LEFT + 1)
`define DSU_CHI_REQ_FLIT_TAGOP_LEFT        (`DSU_CHI_REQ_FLIT_TAGOP_RIGHT + `DSU_CHI_REQ_FLIT_TAGOP_WIDTH - 1)

// TRACETAG
`define DSU_CHI_REQ_FLIT_TRACETAG_RIGHT    (`DSU_CHI_REQ_FLIT_TAGOP_LEFT + 1)
`define DSU_CHI_REQ_FLIT_TRACETAG_LEFT     (`DSU_CHI_REQ_FLIT_TRACETAG_RIGHT + `DSU_CHI_REQ_FLIT_TRACETAG_WIDTH - 1)

//MPAM
`define DSU_CHI_REQ_FLIT_MPAM_RIGHT        (`DSU_CHI_REQ_FLIT_TRACETAG_LEFT + 1)
`define DSU_CHI_REQ_FLIT_MPAM_LEFT         (`DSU_CHI_REQ_FLIT_MPAM_RIGHT + `DSU_CHI_REQ_FLIT_MPAM_WIDTH - 1)

// RSVD
`define DSU_CHI_REQ_FLIT_RSVD_RIGHT        (`DSU_CHI_REQ_FLIT_MPAM_LEFT + 1)
`define DSU_CHI_REQ_FLIT_RSVD_LEFT         (`DSU_CHI_REQ_FLIT_RSVD_RIGHT + `DSU_CHI_REQ_FLIT_RSVD_WIDTH - 1)

// SRCTYPE
`define DSU_CHI_REQ_FLIT_SRCTYPE_RIGHT     (`DSU_CHI_REQ_FLIT_RSVD_LEFT + 1)
`define DSU_CHI_REQ_FLIT_SRCTYPE_LEFT      (`DSU_CHI_REQ_FLIT_SRCTYPE_RIGHT + `DSU_CHI_REQ_FLIT_SRCTYPE_WIDTH - 1)

// LDID
`define DSU_CHI_REQ_FLIT_LDID_RIGHT        (`DSU_CHI_REQ_FLIT_SRCTYPE_LEFT + 1)
`define DSU_CHI_REQ_FLIT_LDID_LEFT         (`DSU_CHI_REQ_FLIT_LDID_RIGHT + `DSU_CHI_REQ_FLIT_LDID_WIDTH - 1)



// RSPQOS
`define DSU_CHI_RSP_FLIT_QOS_RIGHT    0
`define DSU_CHI_RSP_FLIT_QOS_LEFT     (`DSU_CHI_RSP_FLIT_QOS_RIGHT + `DSU_CHI_RSP_FLIT_QOS_WIDTH - 1)

// RSPTGTID
`define DSU_CHI_RSP_FLIT_TGTID_RIGHT      (`DSU_CHI_RSP_FLIT_QOS_LEFT + 1)
`define DSU_CHI_RSP_FLIT_TGTID_LEFT       (`DSU_CHI_RSP_FLIT_TGTID_RIGHT + `DSU_CHI_RSP_FLIT_TGTID_WIDTH - 1)
`define DSU_CHI_RSP_FLIT_DEVICEID_RIGHT   (`DSU_CHI_RSP_FLIT_QOS_LEFT + 1)
`define DSU_CHI_RSP_FLIT_DEVICEID_LEFT    (`DSU_CHI_RSP_FLIT_DEVICEID_RIGHT + `DSU_MXP_DEVICEID_WIDTH_PARAM - 1)
`define DSU_CHI_RSP_FLIT_PORTID_RIGHT     (`DSU_CHI_RSP_FLIT_DEVICEID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_PORTID_LEFT      (`DSU_CHI_RSP_FLIT_PORTID_RIGHT + `DSU_MXP_PORTID_WIDTH_PARAM - 1)
`define DSU_CHI_RSP_FLIT_YID_RIGHT        (`DSU_CHI_RSP_FLIT_PORTID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_YID_LEFT         (`DSU_CHI_RSP_FLIT_YID_RIGHT + `DSU_MXP_YID_WIDTH_PARAM - 1)
`define DSU_CHI_RSP_FLIT_XID_RIGHT        (`DSU_CHI_RSP_FLIT_YID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_XID_LEFT         (`DSU_CHI_RSP_FLIT_XID_RIGHT + `DSU_MXP_XID_WIDTH_PARAM - 1)
`define DSU_CHI_RSP_FLIT_MESHID_RIGHT     (`DSU_CHI_RSP_FLIT_XID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_MESHID_LEFT      (`DSU_CHI_RSP_FLIT_MESHID_RIGHT + `DSU_MXP_MESHID_WIDTH_PARAM - 1)


// RSPSRCID
`define DSU_CHI_RSP_FLIT_SRCID_RIGHT  (`DSU_CHI_RSP_FLIT_TGTID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_SRCID_LEFT   (`DSU_CHI_RSP_FLIT_SRCID_RIGHT + `DSU_CHI_RSP_FLIT_SRCID_WIDTH - 1)

// RSPTXNID
`define DSU_CHI_RSP_FLIT_TXNID_RIGHT  (`DSU_CHI_RSP_FLIT_SRCID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_TXNID_LEFT   (`DSU_CHI_RSP_FLIT_TXNID_RIGHT + `DSU_CHI_RSP_FLIT_TXNID_WIDTH - 1)

// RSPOPCODE
`define DSU_CHI_RSP_FLIT_OPCODE_RIGHT (`DSU_CHI_RSP_FLIT_TXNID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_OPCODE_LEFT  (`DSU_CHI_RSP_FLIT_OPCODE_RIGHT + `DSU_CHI_RSP_FLIT_OPCODE_WIDTH - 1)

// RSPRESPERR
`define DSU_CHI_RSP_FLIT_RESPERR_RIGHT (`DSU_CHI_RSP_FLIT_OPCODE_LEFT + 1)
`define DSU_CHI_RSP_FLIT_RESPERR_LEFT  (`DSU_CHI_RSP_FLIT_RESPERR_RIGHT + `DSU_CHI_RSP_FLIT_RESPERR_WIDTH - 1)

// RSPRESP
`define DSU_CHI_RSP_FLIT_RESP_RIGHT   (`DSU_CHI_RSP_FLIT_RESPERR_LEFT + 1)
`define DSU_CHI_RSP_FLIT_RESP_LEFT    (`DSU_CHI_RSP_FLIT_RESP_RIGHT + `DSU_CHI_RSP_FLIT_RESP_WIDTH - 1)

`define DSU_CHI_RSP_FLIT_RESPSNP_RIGHT   (`DSU_CHI_RSP_FLIT_RESPERR_LEFT + 1)
`define DSU_CHI_RSP_FLIT_RESPSNP_LEFT    (`DSU_CHI_RSP_FLIT_RESPSNP_RIGHT + `DSU_CHI_RSP_FLIT_RESPSNP_WIDTH - 1)  

`define DSU_CHI_RSP_FLIT_RESPPASSDIRTY_RIGHT   (`DSU_CHI_RSP_FLIT_RESPSNP_LEFT + 1)
`define DSU_CHI_RSP_FLIT_RESPPASSDIRTY_LEFT    (`DSU_CHI_RSP_FLIT_RESPPASSDIRTY_RIGHT + `DSU_CHI_RSP_FLIT_RESPPASSDIRTY_WIDTH - 1)  

// RSPFWDSTATE
`define DSU_CHI_RSP_FLIT_FWDSTATE_RIGHT (`DSU_CHI_RSP_FLIT_RESP_LEFT + 1)
`define DSU_CHI_RSP_FLIT_FWDSTATE_LEFT  (`DSU_CHI_RSP_FLIT_FWDSTATE_RIGHT + `DSU_CHI_RSP_FLIT_FWDSTATE_WIDTH - 1)

// RSPCBUSY
`define DSU_CHI_RSP_FLIT_CBUSY_RIGHT   (`DSU_CHI_RSP_FLIT_FWDSTATE_LEFT + 1)
`define DSU_CHI_RSP_FLIT_CBUSY_LEFT    (`DSU_CHI_RSP_FLIT_CBUSY_RIGHT + `DSU_CHI_RSP_FLIT_CBUSY_WIDTH - 1)

// RSPDBID
`define DSU_CHI_RSP_FLIT_DBID_RIGHT   (`DSU_CHI_RSP_FLIT_CBUSY_LEFT + 1)
`define DSU_CHI_RSP_FLIT_DBID_LEFT    (`DSU_CHI_RSP_FLIT_DBID_RIGHT + `DSU_CHI_RSP_FLIT_DBID_WIDTH - 1)

// RSPPCRDTYPE
`define DSU_CHI_RSP_FLIT_PCRDTYPE_RIGHT (`DSU_CHI_RSP_FLIT_DBID_LEFT + 1)
`define DSU_CHI_RSP_FLIT_PCRDTYPE_LEFT  (`DSU_CHI_RSP_FLIT_PCRDTYPE_RIGHT + `DSU_CHI_RSP_FLIT_PCRDTYPE_WIDTH - 1)

// RSPTAGOP
`define DSU_CHI_RSP_FLIT_TAGOP_RIGHT   (`DSU_CHI_RSP_FLIT_PCRDTYPE_LEFT + 1)
`define DSU_CHI_RSP_FLIT_TAGOP_LEFT    (`DSU_CHI_RSP_FLIT_TAGOP_RIGHT + `DSU_CHI_RSP_FLIT_TAGOP_WIDTH - 1)

// RSPTRACETAG
`define DSU_CHI_RSP_FLIT_TRACETAG_RIGHT (`DSU_CHI_RSP_FLIT_TAGOP_LEFT + 1)
`define DSU_CHI_RSP_FLIT_TRACETAG_LEFT  (`DSU_CHI_RSP_FLIT_TRACETAG_RIGHT + `DSU_CHI_RSP_FLIT_TRACETAG_WIDTH - 1)

// RSPDEVEVENT
`define DSU_CHI_RSP_FLIT_DEVEVENT_RIGHT (`DSU_CHI_RSP_FLIT_TRACETAG_LEFT + 1)
`define DSU_CHI_RSP_FLIT_DEVEVENT_LEFT  (`DSU_CHI_RSP_FLIT_DEVEVENT_RIGHT + `DSU_CHI_RSP_FLIT_DEVEVENT_WIDTH - 1)



// DATQOS
`define DSU_CHI_DAT_FLIT_QOS_RIGHT    0
`define DSU_CHI_DAT_FLIT_QOS_LEFT     (`DSU_CHI_DAT_FLIT_QOS_RIGHT + `DSU_CHI_DAT_FLIT_QOS_WIDTH - 1)

// DATTGTID
`define DSU_CHI_DAT_FLIT_TGTID_RIGHT      (`DSU_CHI_DAT_FLIT_QOS_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TGTID_LEFT       (`DSU_CHI_DAT_FLIT_TGTID_RIGHT + `DSU_CHI_DAT_FLIT_TGTID_WIDTH - 1)
`define DSU_CHI_DAT_FLIT_DEVICEID_RIGHT   (`DSU_CHI_DAT_FLIT_QOS_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DEVICEID_LEFT    (`DSU_CHI_DAT_FLIT_DEVICEID_RIGHT + `DSU_MXP_DEVICEID_WIDTH_PARAM - 1)
`define DSU_CHI_DAT_FLIT_PORTID_RIGHT     (`DSU_CHI_DAT_FLIT_DEVICEID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_PORTID_LEFT      (`DSU_CHI_DAT_FLIT_PORTID_RIGHT + `DSU_MXP_PORTID_WIDTH_PARAM - 1)
`define DSU_CHI_DAT_FLIT_YID_RIGHT        (`DSU_CHI_DAT_FLIT_PORTID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_YID_LEFT         (`DSU_CHI_DAT_FLIT_YID_RIGHT + `DSU_MXP_YID_WIDTH_PARAM - 1)
`define DSU_CHI_DAT_FLIT_XID_RIGHT        (`DSU_CHI_DAT_FLIT_YID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_XID_LEFT         (`DSU_CHI_DAT_FLIT_XID_RIGHT + `DSU_MXP_XID_WIDTH_PARAM - 1)
`define DSU_CHI_DAT_FLIT_MESHID_RIGHT     (`DSU_CHI_DAT_FLIT_XID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_MESHID_LEFT      (`DSU_CHI_DAT_FLIT_MESHID_RIGHT + `DSU_MXP_MESHID_WIDTH_PARAM - 1)



// DATSRCID
`define DSU_CHI_DAT_FLIT_SRCID_RIGHT  (`DSU_CHI_DAT_FLIT_TGTID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_SRCID_LEFT   (`DSU_CHI_DAT_FLIT_SRCID_RIGHT + `DSU_CHI_DAT_FLIT_SRCID_WIDTH - 1)

// DATTXNID
`define DSU_CHI_DAT_FLIT_TXNID_RIGHT  (`DSU_CHI_DAT_FLIT_SRCID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TXNID_LEFT   (`DSU_CHI_DAT_FLIT_TXNID_RIGHT + `DSU_CHI_DAT_FLIT_TXNID_WIDTH - 1)

// DATHNID
`define DSU_CHI_DAT_FLIT_HNID_RIGHT   (`DSU_CHI_DAT_FLIT_TXNID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_HNID_LEFT    (`DSU_CHI_DAT_FLIT_HNID_RIGHT + `DSU_CHI_DAT_FLIT_HNID_WIDTH - 1)

// DATOPCODE
`define DSU_CHI_DAT_FLIT_OPCODE_RIGHT (`DSU_CHI_DAT_FLIT_HNID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_OPCODE_LEFT  (`DSU_CHI_DAT_FLIT_OPCODE_RIGHT + `DSU_CHI_DAT_FLIT_OPCODE_WIDTH - 1)

// DATRESPERR
`define DSU_CHI_DAT_FLIT_RESPERR_RIGHT (`DSU_CHI_DAT_FLIT_OPCODE_LEFT + 1)
`define DSU_CHI_DAT_FLIT_RESPERR_LEFT  (`DSU_CHI_DAT_FLIT_RESPERR_RIGHT + `DSU_CHI_DAT_FLIT_RESPERR_WIDTH - 1)

// DATRESP
`define DSU_CHI_DAT_FLIT_RESP_RIGHT   (`DSU_CHI_DAT_FLIT_RESPERR_LEFT + 1)
`define DSU_CHI_DAT_FLIT_RESP_LEFT    (`DSU_CHI_DAT_FLIT_RESP_RIGHT + `DSU_CHI_DAT_FLIT_RESP_WIDTH - 1)

// DATFWDSTATE
`define DSU_CHI_DAT_FLIT_FWDSTATE_RIGHT (`DSU_CHI_DAT_FLIT_RESP_LEFT + 1)
`define DSU_CHI_DAT_FLIT_FWDSTATE_LEFT  (`DSU_CHI_DAT_FLIT_FWDSTATE_RIGHT + `DSU_CHI_DAT_FLIT_FWDSTATE_WIDTH - 1)

// DATCBUSY
`define DSU_CHI_DAT_FLIT_CBUSY_RIGHT   (`DSU_CHI_DAT_FLIT_FWDSTATE_LEFT + 1)
`define DSU_CHI_DAT_FLIT_CBUSY_LEFT    (`DSU_CHI_DAT_FLIT_CBUSY_RIGHT + `DSU_CHI_DAT_FLIT_CBUSY_WIDTH - 1)

// DATDBID
`define DSU_CHI_DAT_FLIT_DBID_RIGHT   (`DSU_CHI_DAT_FLIT_CBUSY_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DBID_LEFT    (`DSU_CHI_DAT_FLIT_DBID_RIGHT + `DSU_CHI_DAT_FLIT_DBID_WIDTH - 1)

// DATCCID
`define DSU_CHI_DAT_FLIT_CCID_RIGHT   (`DSU_CHI_DAT_FLIT_DBID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_CCID_LEFT    (`DSU_CHI_DAT_FLIT_CCID_RIGHT + `DSU_CHI_DAT_FLIT_CCID_WIDTH - 1)

// DATDATAID
`define DSU_CHI_DAT_FLIT_DATAID_RIGHT (`DSU_CHI_DAT_FLIT_CCID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DATAID_LEFT  (`DSU_CHI_DAT_FLIT_DATAID_RIGHT + `DSU_CHI_DAT_FLIT_DATAID_WIDTH - 1)

// DATTAGOP
`define DSU_CHI_DAT_FLIT_TAGOP_RIGHT   (`DSU_CHI_DAT_FLIT_DATAID_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TAGOP_LEFT    (`DSU_CHI_DAT_FLIT_TAGOP_RIGHT + `DSU_CHI_DAT_FLIT_TAGOP_WIDTH - 1)

// DATTAG
`define DSU_CHI_DAT_FLIT_TAG_RIGHT   (`DSU_CHI_DAT_FLIT_TAGOP_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TAG_LEFT    (`DSU_CHI_DAT_FLIT_TAG_RIGHT + `DSU_CHI_DAT_FLIT_TAG_WIDTH - 1)

// DATTU
`define DSU_CHI_DAT_FLIT_TU_RIGHT   (`DSU_CHI_DAT_FLIT_TAG_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TU_LEFT    (`DSU_CHI_DAT_FLIT_TU_RIGHT + `DSU_CHI_DAT_FLIT_TU_WIDTH - 1)

// DATTRACETAG
`define DSU_CHI_DAT_FLIT_TRACETAG_RIGHT (`DSU_CHI_DAT_FLIT_TU_LEFT + 1)
`define DSU_CHI_DAT_FLIT_TRACETAG_LEFT  (`DSU_CHI_DAT_FLIT_TRACETAG_RIGHT + `DSU_CHI_DAT_FLIT_TRACETAG_WIDTH - 1)

// DATRSVD
`define DSU_CHI_DAT_FLIT_RSVD_RIGHT   (`DSU_CHI_DAT_FLIT_TRACETAG_LEFT + 1)
`define DSU_CHI_DAT_FLIT_RSVD_LEFT    (`DSU_CHI_DAT_FLIT_RSVD_RIGHT + `DSU_CHI_DAT_FLIT_RSVD_WIDTH - 1)

// DATBE
`define DSU_CHI_DAT_FLIT_BE_RIGHT     (`DSU_CHI_DAT_FLIT_RSVD_LEFT + 1)
`define DSU_CHI_DAT_FLIT_BE_LEFT      (`DSU_CHI_DAT_FLIT_BE_RIGHT + `DSU_CHI_DAT_FLIT_BE_WIDTH - 1)

// DATDATA
`define DSU_CHI_DAT_FLIT_DATA_RIGHT   (`DSU_CHI_DAT_FLIT_BE_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DATA_LEFT    (`DSU_CHI_DAT_FLIT_DATA_RIGHT + `DSU_CHI_DAT_FLIT_DATA_WIDTH - 1)

// DATDATACHECK
`define DSU_CHI_DAT_FLIT_DATACHECK_RIGHT   (`DSU_CHI_DAT_FLIT_DATA_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DATACHECK_LEFT    (`DSU_CHI_DAT_FLIT_DATACHECK_RIGHT + `DSU_CHI_DAT_FLIT_DATACHECK_WIDTH - 1)

// DATPOISON
`define DSU_CHI_DAT_FLIT_POISON_RIGHT (`DSU_CHI_DAT_FLIT_DATACHECK_LEFT + 1)
`define DSU_CHI_DAT_FLIT_POISON_LEFT  (`DSU_CHI_DAT_FLIT_POISON_RIGHT + `DSU_CHI_DAT_FLIT_POISON_WIDTH - 1)

// DATCHUNKV
`define DSU_CHI_DAT_FLIT_CHUNKV_RIGHT (`DSU_CHI_DAT_FLIT_POISON_LEFT + 1)
`define DSU_CHI_DAT_FLIT_CHUNKV_LEFT  (`DSU_CHI_DAT_FLIT_CHUNKV_RIGHT + `DSU_CHI_DAT_FLIT_CHUNKV_WIDTH - 1)

// DATDEVEVENT
`define DSU_CHI_DAT_FLIT_DEVEVENT_RIGHT (`DSU_CHI_DAT_FLIT_CHUNKV_LEFT + 1)
`define DSU_CHI_DAT_FLIT_DEVEVENT_LEFT  (`DSU_CHI_DAT_FLIT_DEVEVENT_RIGHT + `DSU_CHI_DAT_FLIT_DEVEVENT_WIDTH - 1)



// SNPQOS
`define DSU_CHI_SNP_FLIT_QOS_RIGHT    0
`define DSU_CHI_SNP_FLIT_QOS_LEFT     (`DSU_CHI_SNP_FLIT_QOS_RIGHT + `DSU_CHI_SNP_FLIT_QOS_WIDTH - 1)

// SNPSRCID
`define DSU_CHI_SNP_FLIT_SRCID_RIGHT  (`DSU_CHI_SNP_FLIT_QOS_LEFT + 1)
`define DSU_CHI_SNP_FLIT_SRCID_LEFT   (`DSU_CHI_SNP_FLIT_SRCID_RIGHT + `DSU_CHI_SNP_FLIT_SRCID_WIDTH - 1)

// TSNPXNID
`define DSU_CHI_SNP_FLIT_TXNID_RIGHT  (`DSU_CHI_SNP_FLIT_SRCID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_TXNID_LEFT   (`DSU_CHI_SNP_FLIT_TXNID_RIGHT + `DSU_CHI_SNP_FLIT_TXNID_WIDTH - 1)

// SNPFWDNID
`define DSU_CHI_SNP_FLIT_FWDNID_RIGHT (`DSU_CHI_SNP_FLIT_TXNID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_FWDNID_LEFT  (`DSU_CHI_SNP_FLIT_FWDNID_RIGHT + `DSU_CHI_SNP_FLIT_FWDNID_WIDTH - 1)

// SNPFWDTXNID
`define DSU_CHI_SNP_FLIT_FWDTXNID_RIGHT (`DSU_CHI_SNP_FLIT_FWDNID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_FWDTXNID_LEFT  (`DSU_CHI_SNP_FLIT_FWDTXNID_RIGHT + `DSU_CHI_SNP_FLIT_FWDTXNID_WIDTH - 1)

// SNPOPCODE
`define DSU_CHI_SNP_FLIT_OPCODE_RIGHT (`DSU_CHI_SNP_FLIT_FWDTXNID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_OPCODE_LEFT  (`DSU_CHI_SNP_FLIT_OPCODE_RIGHT + `DSU_CHI_SNP_FLIT_OPCODE_WIDTH - 1)

// SNPADDR
`define DSU_CHI_SNP_FLIT_ADDR_RIGHT   (`DSU_CHI_SNP_FLIT_OPCODE_LEFT + 1)
`define DSU_CHI_SNP_FLIT_ADDR_LEFT    (`DSU_CHI_SNP_FLIT_ADDR_RIGHT + `DSU_CHI_SNP_FLIT_ADDR_WIDTH - 1)

// SNPNS
`define DSU_CHI_SNP_FLIT_NS_RIGHT     (`DSU_CHI_SNP_FLIT_ADDR_LEFT + 1)
`define DSU_CHI_SNP_FLIT_NS_LEFT      (`DSU_CHI_SNP_FLIT_NS_RIGHT + `DSU_CHI_SNP_FLIT_NS_WIDTH - 1)

// SNPDONOTGOTOSD
`define DSU_CHI_SNP_FLIT_DONOTGOTOSD_RIGHT (`DSU_CHI_SNP_FLIT_NS_LEFT + 1)
`define DSU_CHI_SNP_FLIT_DONOTGOTOSD_LEFT  (`DSU_CHI_SNP_FLIT_DONOTGOTOSD_RIGHT + `DSU_CHI_SNP_FLIT_DONOTGOTOSD_WIDTH - 1)

// SNPRETTO_SRC
`define DSU_CHI_SNP_FLIT_RETTO_SRC_RIGHT (`DSU_CHI_SNP_FLIT_DONOTGOTOSD_LEFT + 1)
`define DSU_CHI_SNP_FLIT_RETTO_SRC_LEFT  (`DSU_CHI_SNP_FLIT_RETTO_SRC_RIGHT + `DSU_CHI_SNP_FLIT_RETTO_SRC_WIDTH - 1)

// SNPTRACETAG
`define DSU_CHI_SNP_FLIT_TRACETAG_RIGHT (`DSU_CHI_SNP_FLIT_RETTO_SRC_LEFT + 1)
`define DSU_CHI_SNP_FLIT_TRACETAG_LEFT  (`DSU_CHI_SNP_FLIT_TRACETAG_RIGHT + `DSU_CHI_SNP_FLIT_TRACETAG_WIDTH - 1)

// SNPMPAM
`define DSU_CHI_SNP_FLIT_MPAM_RIGHT (`DSU_CHI_SNP_FLIT_TRACETAG_LEFT + 1)
`define DSU_CHI_SNP_FLIT_MPAM_LEFT  (`DSU_CHI_SNP_FLIT_MPAM_RIGHT + `DSU_CHI_SNP_FLIT_MPAM_WIDTH - 1)

// SNPLDID
`define DSU_CHI_SNP_FLIT_LDID_RIGHT   (`DSU_CHI_SNP_FLIT_MPAM_LEFT + 1)
`define DSU_CHI_SNP_FLIT_LDID_LEFT    (`DSU_CHI_SNP_FLIT_LDID_RIGHT + `DSU_CHI_SNP_FLIT_LDID_WIDTH - 1)

// SNPTGTID
`define DSU_CHI_SNP_FLIT_TGTID_RIGHT      (`DSU_CHI_SNP_FLIT_LDID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_TGTID_LEFT       (`DSU_CHI_SNP_FLIT_TGTID_RIGHT + `DSU_CHI_SNP_FLIT_TGTID_WIDTH - 1)
`define DSU_CHI_SNP_FLIT_DEVICEID_RIGHT   (`DSU_CHI_SNP_FLIT_LDID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_DEVICEID_LEFT    (`DSU_CHI_SNP_FLIT_DEVICEID_RIGHT + `DSU_MXP_DEVICEID_WIDTH_PARAM - 1)
`define DSU_CHI_SNP_FLIT_PORTID_RIGHT     (`DSU_CHI_SNP_FLIT_DEVICEID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_PORTID_LEFT      (`DSU_CHI_SNP_FLIT_PORTID_RIGHT + `DSU_MXP_PORTID_WIDTH_PARAM - 1)
`define DSU_CHI_SNP_FLIT_YID_RIGHT        (`DSU_CHI_SNP_FLIT_PORTID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_YID_LEFT         (`DSU_CHI_SNP_FLIT_YID_RIGHT + `DSU_MXP_YID_WIDTH_PARAM - 1)
`define DSU_CHI_SNP_FLIT_XID_RIGHT        (`DSU_CHI_SNP_FLIT_YID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_XID_LEFT         (`DSU_CHI_SNP_FLIT_XID_RIGHT + `DSU_MXP_XID_WIDTH_PARAM - 1)
`define DSU_CHI_SNP_FLIT_MESHID_RIGHT     (`DSU_CHI_SNP_FLIT_XID_LEFT + 1)
`define DSU_CHI_SNP_FLIT_MESHID_LEFT      (`DSU_CHI_SNP_FLIT_MESHID_RIGHT + `DSU_MXP_MESHID_WIDTH_PARAM - 1)


//Use left and right to indicate range
//REQ
`define DSU_CHI_REQ_FLIT_QOS_RANGE             `DSU_CHI_REQ_FLIT_QOS_LEFT:`DSU_CHI_REQ_FLIT_QOS_RIGHT
`define DSU_CHI_REQ_FLIT_DEVICEID_RANGE        `DSU_CHI_REQ_FLIT_DEVICEID_LEFT:`DSU_CHI_REQ_FLIT_DEVICEID_RIGHT
`define DSU_CHI_REQ_FLIT_PORTID_RANGE          `DSU_CHI_REQ_FLIT_PORTID_LEFT:`DSU_CHI_REQ_FLIT_PORTID_RIGHT
`define DSU_CHI_REQ_FLIT_YID_RANGE             `DSU_CHI_REQ_FLIT_YID_LEFT:`DSU_CHI_REQ_FLIT_YID_RIGHT
`define DSU_CHI_REQ_FLIT_XID_RANGE             `DSU_CHI_REQ_FLIT_XID_LEFT:`DSU_CHI_REQ_FLIT_XID_RIGHT
`define DSU_CHI_REQ_FLIT_MESHID_RANGE          `DSU_CHI_REQ_FLIT_MESHID_LEFT:`DSU_CHI_REQ_FLIT_MESHID_RIGHT
`define DSU_CHI_REQ_FLIT_TGTID_RANGE           `DSU_CHI_REQ_FLIT_TGTID_LEFT:`DSU_CHI_REQ_FLIT_TGTID_RIGHT
`define DSU_CHI_REQ_FLIT_SRCID_RANGE           `DSU_CHI_REQ_FLIT_SRCID_LEFT:`DSU_CHI_REQ_FLIT_SRCID_RIGHT
`define DSU_CHI_REQ_FLIT_TXNID_RANGE           `DSU_CHI_REQ_FLIT_TXNID_LEFT:`DSU_CHI_REQ_FLIT_TXNID_RIGHT
`define DSU_CHI_REQ_FLIT_RNID_RANGE            `DSU_CHI_REQ_FLIT_RNID_LEFT:`DSU_CHI_REQ_FLIT_RNID_RIGHT
`define DSU_CHI_REQ_FLIT_STASHNIDV_RANGE       `DSU_CHI_REQ_FLIT_STASHNIDV_LEFT:`DSU_CHI_REQ_FLIT_STASHNIDV_RIGHT
`define DSU_CHI_REQ_FLIT_STASHLPIDVALID_RANGE  `DSU_CHI_REQ_FLIT_STASHLPIDVALID_LEFT:`DSU_CHI_REQ_FLIT_STASHLPIDVALID_RIGHT
`define DSU_CHI_REQ_FLIT_STASHLPID_RANGE       `DSU_CHI_REQ_FLIT_STASHLPID_LEFT:`DSU_CHI_REQ_FLIT_STASHLPID_RIGHT
`define DSU_CHI_REQ_FLIT_RETURNTXNID_RANGE     `DSU_CHI_REQ_FLIT_RETURNTXNID_LEFT:`DSU_CHI_REQ_FLIT_RETURNTXNID_RIGHT
`define DSU_CHI_REQ_FLIT_OPCODE_RANGE          `DSU_CHI_REQ_FLIT_OPCODE_LEFT:`DSU_CHI_REQ_FLIT_OPCODE_RIGHT
`define DSU_CHI_REQ_FLIT_SIZE_RANGE            `DSU_CHI_REQ_FLIT_SIZE_LEFT:`DSU_CHI_REQ_FLIT_SIZE_RIGHT
`define DSU_CHI_REQ_FLIT_ADDR_RANGE            `DSU_CHI_REQ_FLIT_ADDR_LEFT:`DSU_CHI_REQ_FLIT_ADDR_RIGHT
`define DSU_CHI_REQ_FLIT_NS_RANGE              `DSU_CHI_REQ_FLIT_NS_LEFT:`DSU_CHI_REQ_FLIT_NS_RIGHT
`define DSU_CHI_REQ_FLIT_LS_RANGE              `DSU_CHI_REQ_FLIT_LS_LEFT:`DSU_CHI_REQ_FLIT_LS_RIGHT
`define DSU_CHI_REQ_FLIT_ALLOWRETRY_RANGE      `DSU_CHI_REQ_FLIT_ALLOWRETRY_LEFT:`DSU_CHI_REQ_FLIT_ALLOWRETRY_RIGHT
`define DSU_CHI_REQ_FLIT_ORDER_RANGE           `DSU_CHI_REQ_FLIT_ORDER_LEFT:`DSU_CHI_REQ_FLIT_ORDER_RIGHT
`define DSU_CHI_REQ_FLIT_PCRDTYPE_RANGE        `DSU_CHI_REQ_FLIT_PCRDTYPE_LEFT:`DSU_CHI_REQ_FLIT_PCRDTYPE_RIGHT
`define DSU_CHI_REQ_FLIT_MEMATTR_RANGE         `DSU_CHI_REQ_FLIT_MEMATTR_LEFT:`DSU_CHI_REQ_FLIT_MEMATTR_RIGHT
`define DSU_CHI_REQ_FLIT_MEMATTREWACK_RANGE    `DSU_CHI_REQ_FLIT_MEMATTREWACK_LEFT:`DSU_CHI_REQ_FLIT_MEMATTREWACK_RIGHT             
`define DSU_CHI_REQ_FLIT_MEMATTRCACHE_RANGE    `DSU_CHI_REQ_FLIT_MEMATTRCACHE_LEFT:`DSU_CHI_REQ_FLIT_MEMATTRCACHE_RIGHT             
`define DSU_CHI_REQ_FLIT_MEMATTRALLHINT_RANGE  `DSU_CHI_REQ_FLIT_MEMATTRALLHINT_LEFT:`DSU_CHI_REQ_FLIT_MEMATTRALLHINT_RIGHT        
`define DSU_CHI_REQ_FLIT_MEMATTRDEVICE_RANGE   `DSU_CHI_REQ_FLIT_MEMATTRDEVICE_LEFT:`DSU_CHI_REQ_FLIT_MEMATTRDEVICE_RIGHT           
`define DSU_CHI_REQ_FLIT_SNPATTR_RANGE         `DSU_CHI_REQ_FLIT_SNPATTR_LEFT:`DSU_CHI_REQ_FLIT_SNPATTR_RIGHT
`define DSU_CHI_REQ_FLIT_LPID_RANGE            `DSU_CHI_REQ_FLIT_LPID_LEFT:`DSU_CHI_REQ_FLIT_LPID_RIGHT
`define DSU_CHI_REQ_FLIT_EXCL_RANGE            `DSU_CHI_REQ_FLIT_EXCL_LEFT:`DSU_CHI_REQ_FLIT_EXCL_RIGHT
`define DSU_CHI_REQ_FLIT_EXPCOMPACK_RANGE      `DSU_CHI_REQ_FLIT_EXPCOMPACK_LEFT:`DSU_CHI_REQ_FLIT_EXPCOMPACK_RIGHT
`define DSU_CHI_REQ_FLIT_TAGOP_RANGE           `DSU_CHI_REQ_FLIT_TAGOP_LEFT:`DSU_CHI_REQ_FLIT_TAGOP_RIGHT
`define DSU_CHI_REQ_FLIT_TRACETAG_RANGE        `DSU_CHI_REQ_FLIT_TRACETAG_LEFT:`DSU_CHI_REQ_FLIT_TRACETAG_RIGHT
`define DSU_CHI_REQ_FLIT_MPAM_RANGE            `DSU_CHI_REQ_FLIT_MPAM_LEFT:`DSU_CHI_REQ_FLIT_MPAM_RIGHT
`define DSU_CHI_REQ_FLIT_RSVD_RANGE            `DSU_CHI_REQ_FLIT_RSVD_LEFT:`DSU_CHI_REQ_FLIT_RSVD_RIGHT
`define DSU_CHI_REQ_FLIT_SRCTYPE_RANGE         `DSU_CHI_REQ_FLIT_SRCTYPE_LEFT:`DSU_CHI_REQ_FLIT_SRCTYPE_RIGHT
`define DSU_CHI_REQ_FLIT_LDID_RANGE            `DSU_CHI_REQ_FLIT_LDID_LEFT:`DSU_CHI_REQ_FLIT_LDID_RIGHT

//RSP
`define DSU_CHI_RSP_FLIT_QOS_RANGE           `DSU_CHI_RSP_FLIT_QOS_LEFT:`DSU_CHI_RSP_FLIT_QOS_RIGHT
`define DSU_CHI_RSP_FLIT_DEVICEID_RANGE      `DSU_CHI_RSP_FLIT_DEVICEID_LEFT:`DSU_CHI_RSP_FLIT_DEVICEID_RIGHT
`define DSU_CHI_RSP_FLIT_PORTID_RANGE        `DSU_CHI_RSP_FLIT_PORTID_LEFT:`DSU_CHI_RSP_FLIT_PORTID_RIGHT
`define DSU_CHI_RSP_FLIT_YID_RANGE           `DSU_CHI_RSP_FLIT_YID_LEFT:`DSU_CHI_RSP_FLIT_YID_RIGHT
`define DSU_CHI_RSP_FLIT_XID_RANGE           `DSU_CHI_RSP_FLIT_XID_LEFT:`DSU_CHI_RSP_FLIT_XID_RIGHT
`define DSU_CHI_RSP_FLIT_MESHID_RANGE        `DSU_CHI_RSP_FLIT_MESHID_LEFT:`DSU_CHI_RSP_FLIT_MESHID_RIGHT
`define DSU_CHI_RSP_FLIT_TGTID_RANGE         `DSU_CHI_RSP_FLIT_TGTID_LEFT:`DSU_CHI_RSP_FLIT_TGTID_RIGHT
`define DSU_CHI_RSP_FLIT_SRCID_RANGE         `DSU_CHI_RSP_FLIT_SRCID_LEFT:`DSU_CHI_RSP_FLIT_SRCID_RIGHT
`define DSU_CHI_RSP_FLIT_TXNID_RANGE         `DSU_CHI_RSP_FLIT_TXNID_LEFT:`DSU_CHI_RSP_FLIT_TXNID_RIGHT
`define DSU_CHI_RSP_FLIT_OPCODE_RANGE        `DSU_CHI_RSP_FLIT_OPCODE_LEFT:`DSU_CHI_RSP_FLIT_OPCODE_RIGHT
`define DSU_CHI_RSP_FLIT_RESPERR_RANGE       `DSU_CHI_RSP_FLIT_RESPERR_LEFT:`DSU_CHI_RSP_FLIT_RESPERR_RIGHT
`define DSU_CHI_RSP_FLIT_RESP_RANGE          `DSU_CHI_RSP_FLIT_RESP_LEFT:`DSU_CHI_RSP_FLIT_RESP_RIGHT
`define DSU_CHI_RSP_FLIT_RESPSNP_RANGE       `DSU_CHI_RSP_FLIT_RESPSNP_LEFT:`DSU_CHI_RSP_FLIT_RESPSNP_RIGHT               
`define DSU_CHI_RSP_FLIT_RESPPASSDIRTY_RANGE `DSU_CHI_RSP_FLIT_RESPPASSDIRTY_LEFT:`DSU_CHI_RSP_FLIT_RESPPASSDIRTY_RIGHT   
`define DSU_CHI_RSP_FLIT_FWDSTATE_RANGE      `DSU_CHI_RSP_FLIT_FWDSTATE_LEFT:`DSU_CHI_RSP_FLIT_FWDSTATE_RIGHT
`define DSU_CHI_RSP_FLIT_CBUSY_RANGE         `DSU_CHI_RSP_FLIT_CBUSY_LEFT:`DSU_CHI_RSP_FLIT_CBUSY_RIGHT
`define DSU_CHI_RSP_FLIT_DBID_RANGE          `DSU_CHI_RSP_FLIT_DBID_LEFT:`DSU_CHI_RSP_FLIT_DBID_RIGHT
`define DSU_CHI_RSP_FLIT_PCRDTYPE_RANGE      `DSU_CHI_RSP_FLIT_PCRDTYPE_LEFT:`DSU_CHI_RSP_FLIT_PCRDTYPE_RIGHT
`define DSU_CHI_RSP_FLIT_TAGOP_RANGE         `DSU_CHI_RSP_FLIT_TAGOP_LEFT:`DSU_CHI_RSP_FLIT_TAGOP_RIGHT
`define DSU_CHI_RSP_FLIT_TRACETAG_RANGE      `DSU_CHI_RSP_FLIT_TRACETAG_LEFT:`DSU_CHI_RSP_FLIT_TRACETAG_RIGHT
`define DSU_CHI_RSP_FLIT_DEVEVENT_RANGE      `DSU_CHI_RSP_FLIT_DEVEVENT_LEFT:`DSU_CHI_RSP_FLIT_DEVEVENT_RIGHT

//DAT
`define DSU_CHI_DAT_FLIT_QOS_RANGE           `DSU_CHI_DAT_FLIT_QOS_LEFT:`DSU_CHI_DAT_FLIT_QOS_RIGHT
`define DSU_CHI_DAT_FLIT_DEVICEID_RANGE      `DSU_CHI_DAT_FLIT_DEVICEID_LEFT:`DSU_CHI_DAT_FLIT_DEVICEID_RIGHT
`define DSU_CHI_DAT_FLIT_PORTID_RANGE        `DSU_CHI_DAT_FLIT_PORTID_LEFT:`DSU_CHI_DAT_FLIT_PORTID_RIGHT
`define DSU_CHI_DAT_FLIT_YID_RANGE           `DSU_CHI_DAT_FLIT_YID_LEFT:`DSU_CHI_DAT_FLIT_YID_RIGHT
`define DSU_CHI_DAT_FLIT_XID_RANGE           `DSU_CHI_DAT_FLIT_XID_LEFT:`DSU_CHI_DAT_FLIT_XID_RIGHT
`define DSU_CHI_DAT_FLIT_MESHID_RANGE        `DSU_CHI_DAT_FLIT_MESHID_LEFT:`DSU_CHI_DAT_FLIT_MESHID_RIGHT
`define DSU_CHI_DAT_FLIT_TGTID_RANGE         `DSU_CHI_DAT_FLIT_TGTID_LEFT:`DSU_CHI_DAT_FLIT_TGTID_RIGHT
`define DSU_CHI_DAT_FLIT_SRCID_RANGE         `DSU_CHI_DAT_FLIT_SRCID_LEFT:`DSU_CHI_DAT_FLIT_SRCID_RIGHT
`define DSU_CHI_DAT_FLIT_TXNID_RANGE         `DSU_CHI_DAT_FLIT_TXNID_LEFT:`DSU_CHI_DAT_FLIT_TXNID_RIGHT
`define DSU_CHI_DAT_FLIT_HNID_RANGE          `DSU_CHI_DAT_FLIT_HNID_LEFT:`DSU_CHI_DAT_FLIT_HNID_RIGHT
`define DSU_CHI_DAT_FLIT_OPCODE_RANGE        `DSU_CHI_DAT_FLIT_OPCODE_LEFT:`DSU_CHI_DAT_FLIT_OPCODE_RIGHT
`define DSU_CHI_DAT_FLIT_RESPERR_RANGE       `DSU_CHI_DAT_FLIT_RESPERR_LEFT:`DSU_CHI_DAT_FLIT_RESPERR_RIGHT
`define DSU_CHI_DAT_FLIT_RESP_RANGE          `DSU_CHI_DAT_FLIT_RESP_LEFT:`DSU_CHI_DAT_FLIT_RESP_RIGHT
`define DSU_CHI_DAT_FLIT_FWDSTATE_RANGE      `DSU_CHI_DAT_FLIT_FWDSTATE_LEFT:`DSU_CHI_DAT_FLIT_FWDSTATE_RIGHT
`define DSU_CHI_DAT_FLIT_CBUSY_RANGE         `DSU_CHI_DAT_FLIT_CBUSY_LEFT:`DSU_CHI_DAT_FLIT_CBUSY_RIGHT
`define DSU_CHI_DAT_FLIT_DBID_RANGE          `DSU_CHI_DAT_FLIT_DBID_LEFT:`DSU_CHI_DAT_FLIT_DBID_RIGHT
`define DSU_CHI_DAT_FLIT_CCID_RANGE          `DSU_CHI_DAT_FLIT_CCID_LEFT:`DSU_CHI_DAT_FLIT_CCID_RIGHT
`define DSU_CHI_DAT_FLIT_DATAID_RANGE        `DSU_CHI_DAT_FLIT_DATAID_LEFT:`DSU_CHI_DAT_FLIT_DATAID_RIGHT
`define DSU_CHI_DAT_FLIT_TAGOP_RANGE         `DSU_CHI_DAT_FLIT_TAGOP_LEFT:`DSU_CHI_DAT_FLIT_TAGOP_RIGHT
`define DSU_CHI_DAT_FLIT_TAG_RANGE           `DSU_CHI_DAT_FLIT_TAG_LEFT:`DSU_CHI_DAT_FLIT_TAG_RIGHT
`define DSU_CHI_DAT_FLIT_TU_RANGE            `DSU_CHI_DAT_FLIT_TU_LEFT:`DSU_CHI_DAT_FLIT_TU_RIGHT
`define DSU_CHI_DAT_FLIT_TRACETAG_RANGE      `DSU_CHI_DAT_FLIT_TRACETAG_LEFT:`DSU_CHI_DAT_FLIT_TRACETAG_RIGHT
`define DSU_CHI_DAT_FLIT_RSVD_RANGE          `DSU_CHI_DAT_FLIT_RSVD_LEFT:`DSU_CHI_DAT_FLIT_RSVD_RIGHT
`define DSU_CHI_DAT_FLIT_BE_RANGE            `DSU_CHI_DAT_FLIT_BE_LEFT:`DSU_CHI_DAT_FLIT_BE_RIGHT
`define DSU_CHI_DAT_FLIT_DATA_RANGE          `DSU_CHI_DAT_FLIT_DATA_LEFT:`DSU_CHI_DAT_FLIT_DATA_RIGHT
`define DSU_CHI_DAT_FLIT_DATACHECK_RANGE     `DSU_CHI_DAT_FLIT_DATACHECK_LEFT:`DSU_CHI_DAT_FLIT_DATACHECK_RIGHT
`define DSU_CHI_DAT_FLIT_POISON_RANGE        `DSU_CHI_DAT_FLIT_POISON_LEFT:`DSU_CHI_DAT_FLIT_POISON_RIGHT
`define DSU_CHI_DAT_FLIT_CHUNKV_RANGE        `DSU_CHI_DAT_FLIT_CHUNKV_LEFT:`DSU_CHI_DAT_FLIT_CHUNKV_RIGHT
`define DSU_CHI_DAT_FLIT_DEVEVENT_RANGE      `DSU_CHI_DAT_FLIT_DEVEVENT_LEFT:`DSU_CHI_DAT_FLIT_DEVEVENT_RIGHT

//SNP
`define DSU_CHI_SNP_FLIT_QOS_RANGE           `DSU_CHI_SNP_FLIT_QOS_LEFT:`DSU_CHI_SNP_FLIT_QOS_RIGHT
`define DSU_CHI_SNP_FLIT_SRCID_RANGE         `DSU_CHI_SNP_FLIT_SRCID_LEFT:`DSU_CHI_SNP_FLIT_SRCID_RIGHT
`define DSU_CHI_SNP_FLIT_TXNID_RANGE         `DSU_CHI_SNP_FLIT_TXNID_LEFT:`DSU_CHI_SNP_FLIT_TXNID_RIGHT
`define DSU_CHI_SNP_FLIT_FWDNID_RANGE        `DSU_CHI_SNP_FLIT_FWDNID_LEFT:`DSU_CHI_SNP_FLIT_FWDNID_RIGHT
`define DSU_CHI_SNP_FLIT_FWDTXNID_RANGE      `DSU_CHI_SNP_FLIT_FWDTXNID_LEFT:`DSU_CHI_SNP_FLIT_FWDTXNID_RIGHT
`define DSU_CHI_SNP_FLIT_OPCODE_RANGE        `DSU_CHI_SNP_FLIT_OPCODE_LEFT:`DSU_CHI_SNP_FLIT_OPCODE_RIGHT
`define DSU_CHI_SNP_FLIT_ADDR_RANGE          `DSU_CHI_SNP_FLIT_ADDR_LEFT:`DSU_CHI_SNP_FLIT_ADDR_RIGHT
`define DSU_CHI_SNP_FLIT_NS_RANGE            `DSU_CHI_SNP_FLIT_NS_LEFT:`DSU_CHI_SNP_FLIT_NS_RIGHT
`define DSU_CHI_SNP_FLIT_DONOTGOTOSD_RANGE   `DSU_CHI_SNP_FLIT_DONOTGOTOSD_LEFT:`DSU_CHI_SNP_FLIT_DONOTGOTOSD_RIGHT
`define DSU_CHI_SNP_FLIT_RETTO_SRC_RANGE     `DSU_CHI_SNP_FLIT_RETTO_SRC_LEFT:`DSU_CHI_SNP_FLIT_RETTO_SRC_RIGHT
`define DSU_CHI_SNP_FLIT_TRACETAG_RANGE      `DSU_CHI_SNP_FLIT_TRACETAG_LEFT:`DSU_CHI_SNP_FLIT_TRACETAG_RIGHT
`define DSU_CHI_SNP_FLIT_MPAM_RANGE          `DSU_CHI_SNP_FLIT_MPAM_LEFT:`DSU_CHI_SNP_FLIT_MPAM_RIGHT
`define DSU_CHI_SNP_FLIT_LDID_RANGE          `DSU_CHI_SNP_FLIT_LDID_LEFT:`DSU_CHI_SNP_FLIT_LDID_RIGHT
`define DSU_CHI_SNP_FLIT_DEVICEID_RANGE      `DSU_CHI_SNP_FLIT_DEVICEID_LEFT:`DSU_CHI_SNP_FLIT_DEVICEID_RIGHT
`define DSU_CHI_SNP_FLIT_PORTID_RANGE        `DSU_CHI_SNP_FLIT_PORTID_LEFT:`DSU_CHI_SNP_FLIT_PORTID_RIGHT
`define DSU_CHI_SNP_FLIT_YID_RANGE           `DSU_CHI_SNP_FLIT_YID_LEFT:`DSU_CHI_SNP_FLIT_YID_RIGHT
`define DSU_CHI_SNP_FLIT_XID_RANGE           `DSU_CHI_SNP_FLIT_XID_LEFT:`DSU_CHI_SNP_FLIT_XID_RIGHT
`define DSU_CHI_SNP_FLIT_MESHID_RANGE        `DSU_CHI_SNP_FLIT_MESHID_LEFT:`DSU_CHI_SNP_FLIT_MESHID_RIGHT
`define DSU_CHI_SNP_FLIT_TGTID_RANGE         `DSU_CHI_SNP_FLIT_TGTID_LEFT:`DSU_CHI_SNP_FLIT_TGTID_RIGHT


//MEMATTR
`define DSU_CHI_MEMATTR_ALLOCATE_RANGE         3
`define DSU_CHI_MEMATTR_CACHEABLE_RANGE        2
`define DSU_CHI_MEMATTR_DEVICE_RANGE           1
`define DSU_CHI_MEMATTR_EARLYWRACK_RANGE       0

//opcode
//TXDAT opcode
`define DSU_CHI_DAT_OP_DATLCRDRETURN           4'h0
`define DSU_CHI_DAT_OP_SNPRESPDATA             4'h1
`define DSU_CHI_DAT_OP_CBWRDATA                4'h2
`define DSU_CHI_DAT_OP_NONCBWRDATA             4'h3
`define DSU_CHI_DAT_OP_COMPDATA                4'h4
`define DSU_CHI_DAT_OP_SNPRSPDATAPTL           4'h5
`define DSU_CHI_DAT_OP_SNPRESPDATAFWDED        4'h6
`define DSU_CHI_DAT_OP_WRITEDATACANCEL         4'h7
`define DSU_CHI_DAT_OP_DATASEPRESP             4'hb
`define DSU_CHI_DAT_OP_NCBWRDATACOMPACK        4'hc
//TXSNP opcode
`define DSU_CHI_SNP_OP_SNPLCRDRETURN           5'h00
`define DSU_CHI_SNP_OP_SNPSHARED               5'h01
`define DSU_CHI_SNP_OP_SNPCLEAN                5'h02
`define DSU_CHI_SNP_OP_SNPONCE                 5'h03
`define DSU_CHI_SNP_OP_SNPNOTSHAREDDIRTY       5'h04
`define DSU_CHI_SNP_OP_SNPUNIQUESTASH          5'h05
`define DSU_CHI_SNP_OP_SNPMAKEINVALIDSTASH     5'h06
`define DSU_CHI_SNP_OP_SNPUNIQUE               5'h07
`define DSU_CHI_SNP_OP_SNPCLEANSHARED          5'h08
`define DSU_CHI_SNP_OP_SNPCLEANINVALID         5'h09
`define DSU_CHI_SNP_OP_SNPMAKEINVALID          5'h0a
`define DSU_CHI_SNP_OP_SNPSTASHUNIQUE          5'h0b
`define DSU_CHI_SNP_OP_SNPSTASHSHARED          5'h0c
`define DSU_CHI_SNP_OP_SNPDVMOP                5'h0d
`define DSU_CHI_SNP_OP_SNPQUERY                5'h10
`define DSU_CHI_SNP_OP_SNPSHAREDFWD            5'h11
`define DSU_CHI_SNP_OP_SNPCLEANFWD             5'h12
`define DSU_CHI_SNP_OP_SNPONCEFWD              5'h13
`define DSU_CHI_SNP_OP_SNPNOTSHAREDDIRTYFWD    5'h14
`define DSU_CHI_SNP_OP_SNPPREFERUNIQUE         5'h15
`define DSU_CHI_SNP_OP_SNPPREFERUNIQUEFWD      5'h16
`define DSU_CHI_SNP_OP_SNPUNIQUEFWD            5'h17
//TXRSP opcode
`define DSU_CHI_RSP_OP_RSPLCRDRETURN           5'h00
`define DSU_CHI_RSP_OP_SNPRESP                 5'h01
`define DSU_CHI_RSP_OP_COMPACK                 5'h02
`define DSU_CHI_RSP_OP_RETRYACK                5'h03
`define DSU_CHI_RSP_OP_COMP                    5'h04
`define DSU_CHI_RSP_OP_COMPDBIDRESP            5'h05
`define DSU_CHI_RSP_OP_DBIDRESP                5'h06
`define DSU_CHI_RSP_OP_CRDGNT                  5'h07
`define DSU_CHI_RSP_OP_READRECEIPT             5'h08
`define DSU_CHI_RSP_OP_SNPRESPFWDED            5'h09
`define DSU_CHI_RSP_OP_TAGMATCH                5'h0a
`define DSU_CHI_RSP_OP_RESPSEPDATA             5'h0b
`define DSU_CHI_RSP_OP_PERSIST                 5'h0c
`define DSU_CHI_RSP_OP_COMPPERSIST             5'h0d
`define DSU_CHI_RSP_OP_DBIDRESPORD             5'h0e
`define DSU_CHI_RSP_OP_STASHDONE               5'h10
`define DSU_CHI_RSP_OP_COMPSTASHDONE           5'h11
`define DSU_CHI_RSP_OP_COMPCMP                 5'h14
//TXREQ opcode
`define DSU_CHI_REQ_OP_REQLCRDRETURN                  7'h00
`define DSU_CHI_REQ_OP_READSHARED                     7'h01
`define DSU_CHI_REQ_OP_READCLEAN                      7'h02
`define DSU_CHI_REQ_OP_READONCE                       7'h03
`define DSU_CHI_REQ_OP_READNOSNP                      7'h04
`define DSU_CHI_REQ_OP_PCRDRETURN                     7'h05
`define DSU_CHI_REQ_OP_READUNIQUE                     7'h07
`define DSU_CHI_REQ_OP_CLEANSHARED                    7'h08
`define DSU_CHI_REQ_OP_CLEANINVALID                   7'h09
`define DSU_CHI_REQ_OP_MAKEINVALID                    7'h0a
`define DSU_CHI_REQ_OP_CLEANUNIQUE                    7'h0b
`define DSU_CHI_REQ_OP_MAKEUNIQUE                     7'h0c
`define DSU_CHI_REQ_OP_EVICT                          7'h0d
`define DSU_CHI_REQ_OP_EOBARRIER                      7'h0e
`define DSU_CHI_REQ_OP_ECBARRIER                      7'h0f
`define DSU_CHI_REQ_OP_READNOSNPSEP                   7'h11
`define DSU_CHI_REQ_OP_CLEANSHAREDPERSISTSEP          7'h13
`define DSU_CHI_REQ_OP_DVMOP                          7'h14
`define DSU_CHI_REQ_OP_EVICTDATAUC                    7'h15
`define DSU_CHI_REQ_OP_WRITEEVICTFULL                 7'h15
`define DSU_CHI_REQ_OP_WRITECLEANFULL                 7'h17
`define DSU_CHI_REQ_OP_WRITEUNIQUEPTL                 7'h18
`define DSU_CHI_REQ_OP_WRITEUNIQUEFULL                7'h19
`define DSU_CHI_REQ_OP_WRITEBACKPTL                   7'h1a
`define DSU_CHI_REQ_OP_WRITEBACKFULL                  7'h1b
`define DSU_CHI_REQ_OP_WRITENOSNPPTL                  7'h1c
`define DSU_CHI_REQ_OP_WRITENOSNPFULL                 7'h1d
`define DSU_CHI_REQ_OP_WRITEUNIQUEFULLSTASH           7'h20
`define DSU_CHI_REQ_OP_WRITEUNIQUEPTLSTASH            7'h21
`define DSU_CHI_REQ_OP_STASHONCESHARED                7'h22
`define DSU_CHI_REQ_OP_STASHONCEUNIQUE                7'h23
`define DSU_CHI_REQ_OP_READONCECLEANINVALID           7'h24
`define DSU_CHI_REQ_OP_READONCEMAKEINVALID            7'h25
`define DSU_CHI_REQ_OP_READNOTSHAREDDIRTY             7'h26
`define DSU_CHI_REQ_OP_CLEANSHAREDPERSIST             7'h27
`define DSU_CHI_REQ_OP_PREFETCHTGT                    7'h3a
`define DSU_CHI_REQ_OP_MAKEREADUNIQUE                 7'h41
`define DSU_CHI_REQ_OP_WRITEEVICTOREVICT              7'h42
`define DSU_CHI_REQ_OP_WRITEUNIQUEZERO                7'h43
`define DSU_CHI_REQ_OP_WRITENOSNPZERO                 7'h44
`define DSU_CHI_REQ_OP_STASHONCESEPSHARED             7'h47
`define DSU_CHI_REQ_OP_STASHONCESEPUNIQUE             7'h48
`define DSU_CHI_REQ_OP_READPREFERUNIQUE               7'h4c
`define DSU_CHI_REQ_OP_WRITENOSNPFULLCLEANSH          7'h50
`define DSU_CHI_REQ_OP_WRITENOSNPFULLCLEANINV         7'h51
`define DSU_CHI_REQ_OP_WRITENOSNPFULLCLEANSHPERSEP    7'h52
`define DSU_CHI_REQ_OP_WRITEUNIQUEFULLCLEANSH         7'h54
`define DSU_CHI_REQ_OP_WRITEUNIQUEFULLCLEANSHPERSEP   7'h56
`define DSU_CHI_REQ_OP_WRITEBACKFULLCLEANSH           7'h58
`define DSU_CHI_REQ_OP_WRITEBACKFULLCLEANINV          7'h59
`define DSU_CHI_REQ_OP_WRITEBACKFULLCLEANSHPERSEP     7'h5a
`define DSU_CHI_REQ_OP_WRITECLEANFULLCLEANSH          7'h5c
`define DSU_CHI_REQ_OP_WRITECLEANFULLCLEANSHPERSEP    7'h5e
`define DSU_CHI_REQ_OP_WRITENOSNPPTLCLEANSH           7'h60
`define DSU_CHI_REQ_OP_WRITENOSNPPTLCLEANINV          7'h61
`define DSU_CHI_REQ_OP_WRITENOSNPPTLCLEANSHPERSEP     7'h62
`define DSU_CHI_REQ_OP_WRITEUNIQUEPTLCLEANSH          7'h64
`define DSU_CHI_REQ_OP_WRITEUNIQUEPTLCLEANSHPERSEP    7'h66

//DAIA SIZE
`define DSU_CHI_DAT_DEFAULT_SIZE               3'b110
`define DSU_CHI_DAT_SIZE1B                     3'h0
`define DSU_CHI_DAT_SIZE2B                     3'h1
`define DSU_CHI_DAT_SIZE4B                     3'h2
`define DSU_CHI_DAT_SIZE8B                     3'h3
`define DSU_CHI_DAT_SIZE16B                    3'h4
`define DSU_CHI_DAT_SIZE32B                    3'h5
`define DSU_CHI_DAT_SIZE64B                    3'h6

